blah

vCLK CLK 0 pulse(0 2.5V 0.5ns 150ps 150ps 0.350ns 1ns )
vVDD VDD! 0 DC 2.5V
vGND GND! 0 DC 0
.OPTION list post=2   
.tran 0.01p 24n
.measure tran avgpwr AVG power from=0ns to=24ns
 
.lib 'models25.txt' TT
   
   
C44 0 2  41.904E-18 M=1.0 
C45 0 1  26.1900000000002E-18 M=1.0 
C46 0 Q3N  32.1264E-18 M=1.0 
C47 0 Q1DOUBLEINV  41.904E-18 M=1.0 
C48 0 XOROUT  29.3328E-18 M=1.0 
C49 CKON 0  226.2816E-18 M=1.0 
C50 VDD! 2  36.3168E-18 M=1.0 
C51 VDD! 1  40.8564E-18 M=1.0 
C52 VDD! Q3N  29.3328E-18 M=1.0 
C53 VDD! XOROUT  41.904E-18 M=1.0 
C54 VDD! CKON  173.2032E-18 M=1.0 
C55 Q2N 0  32.1264E-18 M=1.0 
C56 Q2N VDD!  29.3328E-18 M=1.0 
C57 Q5 0  32.1264E-18 M=1.0 
C58 Q5 VDD!  29.3328E-18 M=1.0 
C59 Q4 0  32.1264E-18 M=1.0 
C60 Q4 VDD!  29.3328E-18 M=1.0 
C61 Q3 0  67.0464E-18 M=1.0 
C62 Q3 VDD!  61.4592E-18 M=1.0 
C63 Q2 0  32.1264E-18 M=1.0 
C64 Q2 VDD!  29.3328000000001E-18 M=1.0 
C65 Q1 0  34.92E-18 M=1.0 
C66 Q1 VDD!  32.1264E-18 M=1.0 
C67 Q1N 0  32.1264000000001E-18 M=1.0 
C68 Q1N VDD!  29.3328000000001E-18 M=1.0 
C69 OUT 0  26.5391999999999E-18 M=1.0 
C70 OUT VDD!  48.8879999999999E-18 M=1.0 
C71 CLK 0  47.4912E-18 M=1.0 
C72 CLK VDD!  78.2208E-18 M=1.0 
C73 CKO 0  262.9476E-18 M=1.0 
C74 CKO VDD!  197.9964E-18 M=1.0 
C75 Q1INV 0  34.92E-18 M=1.0 
C76 Q1INV VDD!  67.0464E-18 M=1.0 
C77 XORINV 0  33.5232E-18 M=1.0 
C78 XORINV VDD!  27.936E-18 M=1.0 
C79 Q3INV 0  34.9199999999999E-18 M=1.0 
C80 Q3INV VDD!  33.5232E-18 M=1.0 
C81 Q5N 0  32.1264E-18 M=1.0 
C82 Q5N VDD!  29.3328E-18 M=1.0 
C83 Q4N 0  32.1264000000001E-18 M=1.0 
C84 Q4N VDD!  29.3328E-18 M=1.0 
C85 0 2  38.0448E-18 M=1.0 
C86 0 1  83.9232E-18 M=1.0 
C87 0 Q3N  90.96E-18 M=1.0 
C88 0 Q1DOUBLEINV  365.2416E-18 M=1.0 
C89 0 XOROUT  133.3824E-18 M=1.0 
C90 CKON 0  290.2848E-18 M=1.0 
C91 VDD! 2  45.2064E-18 M=1.0 
C92 VDD! 1  94.9392E-18 M=1.0 
C93 VDD! Q3N  92.0304E-18 M=1.0 
C94 VDD! Q1DOUBLEINV  51.2496E-18 M=1.0 
C95 VDD! XOROUT  144.1488E-18 M=1.0 
C96 VDD! CKON  267.336E-18 M=1.0 
C97 Q2N 0  90.96E-18 M=1.0 
C98 Q2N VDD!  92.0304E-18 M=1.0 
C99 Q5 0  90.96E-18 M=1.0 
C100 Q5 VDD!  92.0304E-18 M=1.0 
C101 Q4 0  91.4952E-18 M=1.0 
C102 Q4 VDD!  91.4952E-18 M=1.0 
C103 Q3 0  438.3888E-18 M=1.0 
C104 Q3 VDD!  318.4128E-18 M=1.0 
C105 Q2 0  90.96E-18 M=1.0 
C106 Q2 VDD!  92.0304E-18 M=1.0 
C107 Q1 0  102.5472E-18 M=1.0 
C108 Q1 VDD!  211.2912E-18 M=1.0 
C109 Q1N 0  90.96E-18 M=1.0 
C110 Q1N VDD!  92.0304E-18 M=1.0 
C111 OUT VDD!  38.0448E-18 M=1.0 
C112 CKO 0  428.58E-18 M=1.0 
C113 CKO VDD!  196.8264E-18 M=1.0 
C114 Q1INV 0  148.3008E-18 M=1.0 
C115 Q1INV VDD!  521.7264E-18 M=1.0 
C116 XORINV 0  472.404E-18 M=1.0 
C117 XORINV VDD!  110.8152E-18 M=1.0 
C118 Q3INV 0  213.4992E-18 M=1.0 
C119 Q3INV VDD!  200.1624E-18 M=1.0 
C120 Q3INV Q1INV  42.9072E-18 M=1.0 
C121 Q5N 0  91.4952E-18 M=1.0 
C122 Q5N VDD!  91.4952E-18 M=1.0 
C123 Q4N 0  90.96E-18 M=1.0 
C124 Q4N VDD!  92.0304E-18 M=1.0 
C125 0 2  104.0472E-18 M=1.0 
C126 0 Q3N  146.3424E-18 M=1.0 
C127 0 XOROUT  711.0936E-18 M=1.0 
C128 CKON Q3N  252.9912E-18 M=1.0 
C129 CKON 0  1.8614088E-15 M=1.0 
C130 VDD! 2  95.7528E-18 M=1.0 
C131 VDD! Q3N  146.4864E-18 M=1.0 
C132 VDD! XOROUT  435.5808E-18 M=1.0 
C133 VDD! CKON  2.1848232E-15 M=1.0 
C134 Q2N 0  146.3424E-18 M=1.0 
C135 Q2N CKON  252.9912E-18 M=1.0 
C136 Q2N VDD!  146.4864E-18 M=1.0 
C137 Q5 0  146.3424E-18 M=1.0 
C138 Q5 CKON  238.9128E-18 M=1.0 
C139 Q5 VDD!  146.4864E-18 M=1.0 
C140 Q4 0  146.3424E-18 M=1.0 
C141 Q4 CKON  234.5376E-18 M=1.0 
C142 Q4 VDD!  146.4864E-18 M=1.0 
C143 Q3 XOROUT  131.544E-18 M=1.0 
C144 Q3 0  146.3424E-18 M=1.0 
C145 Q3 CKON  238.9128E-18 M=1.0 
C146 Q3 VDD!  146.4864E-18 M=1.0 
C147 Q2 0  146.3424E-18 M=1.0 
C148 Q2 CKON  238.9128E-18 M=1.0 
C149 Q2 VDD!  146.4864E-18 M=1.0 
C150 Q1 0  146.3424E-18 M=1.0 
C151 Q1 VDD!  146.364E-18 M=1.0 
C152 Q1N 2  120.8448E-18 M=1.0 
C153 Q1N 0  146.3424E-18 M=1.0 
C154 Q1N CKON  51.5184E-18 M=1.0 
C155 Q1N VDD!  146.4864E-18 M=1.0 
C156 OUT 0  51.8688E-18 M=1.0 
C157 OUT CKON  51.8688E-18 M=1.0 
C158 OUT VDD!  51.8688E-18 M=1.0 
C159 CKO 0  259.344E-18 M=1.0 
C160 CKO VDD!  259.344E-18 M=1.0 
C161 Q1INV Q1DOUBLEINV  79.6752E-18 M=1.0 
C162 Q1INV XOROUT  133.0272E-18 M=1.0 
C163 Q1INV 0  166.8768E-18 M=1.0 
C164 Q1INV VDD!  169.3536E-18 M=1.0 
C165 Q3INV XOROUT  320.5344E-18 M=1.0 
C166 Q3INV 0  118.4832E-18 M=1.0 
C167 Q3INV VDD!  118.4832E-18 M=1.0 
C168 Q5N 0  146.3424E-18 M=1.0 
C169 Q5N CKON  247.5504E-18 M=1.0 
C170 Q5N VDD!  146.4864E-18 M=1.0 
C171 Q4N 0  146.3424E-18 M=1.0 
C172 Q4N CKON  252.9912E-18 M=1.0 
C173 Q4N VDD!  146.4864E-18 M=1.0 
C174 0 2  336.9168E-18 M=1.0 
C175 0 1  265.7304E-18 M=1.0 
C176 CKON 1  90.648E-18 M=1.0 
C177 CKON 0  1.3476672E-15 M=1.0 
C178 VDD! 2  298.9152E-18 M=1.0 
C179 VDD! 1  269.3808E-18 M=1.0 
C180 VDD! CKON  1.3068792E-15 M=1.0 
C181 OUT 0  63.0072E-18 M=1.0 
C182 OUT VDD!  210.6936E-18 M=1.0 
C183 CLK 1  73.728E-18 M=1.0 
C184 CKO 1  90.648E-18 M=1.0 
C185 XORINV OUT  90.648E-18 M=1.0 
C186 CKO 2  108.048E-18 M=1.0 
C187 CKO 0  1.6200552E-15 M=1.0 
C188 CKO CKON  2.125308E-15 M=1.0 
C189 CKO VDD!  1.308792E-15 M=1.0 
C190 CKO Q5  21.1392E-18 M=1.0 
C191 CKO Q3  21.1392E-18 M=1.0 
C192 CKO Q2  21.1392E-18 M=1.0 
C193 CKO Q1N  70.776E-18 M=1.0 
C194 CKO OUT  104.5536E-18 M=1.0 
C195 0 1  94.0464E-18 M=1.0 
C196 CKON 0  94.1904E-18 M=1.0 
C197 VDD! 1  80.28E-18 M=1.0 
C198 VDD! 0  44.58E-18 M=1.0 
C199 VDD! CKON  94.9824E-18 M=1.0 
C200 Q5 0  112.9752E-18 M=1.0 
C201 CLK 0  92.3616E-18 M=1.0 
C202 CLK VDD!  92.3616E-18 M=1.0 
C203 CKO 0  761.1552E-18 M=1.0 
C204 CKO VDD!  80.7984E-18 M=1.0 
C205 XORINV 0  41.5296E-18 M=1.0 
M206 VDD! XORINV OUT VDD!  pmos  L=239.99999143598E-9 
+W=2.88000001091859E-6 AD=1.72800001304457E-12 AS=1.72800001304457E-12 
+PD=4.08000005336362E-6 PS=4.08000005336362E-6 M=1 
M207 VDD! XOROUT XORINV VDD!  pmos  L=239.99999143598E-9 
+W=1.4400000054593E-6 AD=864.000006522286E-15 AS=864.000006522286E-15 
+PD=2.64000004790432E-6 PS=2.64000004790432E-6 M=1 
M208 VDD! Q1 Q1INV VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=432.000003261143E-15 PD=1.91999993148784E-6 
+PS=1.91999993148784E-6 M=1 
M209 VDD! Q3N 17 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M210 17 CKON Q3 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M211 VDD! OUT 43 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M212 VDD! Q3 16 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M213 43 CKO Q5N VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M214 16 CKO Q2N VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M215 VDD! Q5N 21 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M216 VDD! Q2N 15 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M217 21 CKON Q5 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M218 15 CKON Q2 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M219 VDD! Q5 20 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M220 VDD! Q2 14 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M221 20 CKO Q4N VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M222 14 CKO Q1N VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M223 VDD! Q4N 19 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M224 VDD! Q1N 13 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M225 19 CKON Q4 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M226 13 2 Q1 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M227 VDD! Q4 18 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M228 18 CKO Q3N VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M229 Q1DOUBLEINV Q1INV VDD! VDD!  pmos  L=239.99999143598E-9 
+W=720.000002729648E-9 AD=432.000003261143E-15 AS=432.000003261143E-15 
+PD=1.91999993148784E-6 PS=1.91999993148784E-6 M=1 
M230 VDD! Q3 Q3INV VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=432.000003261143E-15 PD=1.91999993148784E-6 
+PS=1.91999993148784E-6 M=1 
M231 Q3INV Q1INV XOROUT VDD!  pmos  L=239.99999143598E-9 
+W=720.000002729648E-9 AD=432.000003261143E-15 AS=432.000003261143E-15 
+PD=1.91999993148784E-6 PS=1.91999993148784E-6 M=1 
M232 Q1INV Q3INV XOROUT VDD!  pmos  L=239.99999143598E-9 
+W=720.000002729648E-9 AD=432.000003261143E-15 AS=432.000003261143E-15 
+PD=1.91999993148784E-6 PS=1.91999993148784E-6 M=1 
M233 CKO 1 VDD! VDD!  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M234 1 CLK VDD! VDD!  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=388.799994803513E-15 PD=2.27999998969608E-6 
+PS=720.000002729648E-9 M=1 
M235 VDD! CLK CKON VDD!  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=388.799994803513E-15 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M236 CKON CKO VDD! VDD!  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=388.799994803513E-15 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M237 VDD! CKON CKO VDD!  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=388.799994803513E-15 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M238 0 XORINV OUT 0  nmos  L=239.99999143598E-9 W=1.4400000054593E-6 
+AD=864.000006522286E-15 AS=864.000006522286E-15 PD=2.64000004790432E-6 
+PS=2.64000004790432E-6 M=1 
M239 0 XOROUT XORINV 0  nmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=432.000003261143E-15 PD=1.91999993148784E-6 
+PS=1.91999993148784E-6 M=1 
M240 0 Q1 Q1INV 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M241 7 CKO Q3 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M242 0 OUT 12 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M243 0 Q3 6 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M244 12 CKON Q5N 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M245 6 CKON Q2N 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M246 0 Q5N 11 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M247 0 Q2N 5 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M248 11 CKO Q5 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M249 5 CKO Q2 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M250 0 Q5 10 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M251 0 Q2 4 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M252 10 CKON Q4N 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M253 4 2 Q1N 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M254 0 Q4N 9 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M255 0 Q1N 3 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M256 9 CKO Q4 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M257 3 CKO Q1 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M258 0 Q4 8 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M259 8 CKON Q3N 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M260 0 Q3N 7 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M261 Q1DOUBLEINV Q1INV 0 0  nmos  L=239.99999143598E-9 
+W=360.000001364824E-9 AD=273.599990319867E-15 AS=273.599990319867E-15 
+PD=1.7999999499807E-6 PS=1.7999999499807E-6 M=1 
M262 Q3INV Q1DOUBLEINV XOROUT 0  nmos  L=239.99999143598E-9 
+W=360.000001364824E-9 AD=273.599990319867E-15 AS=273.599990319867E-15 
+PD=1.7999999499807E-6 PS=1.7999999499807E-6 M=1 
M263 Q1DOUBLEINV Q3INV XOROUT 0  nmos  L=239.99999143598E-9 
+W=360.000001364824E-9 AD=273.599990319867E-15 AS=273.599990319867E-15 
+PD=1.7999999499807E-6 PS=1.7999999499807E-6 M=1 
M264 0 Q3 Q3INV 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M265 1 CLK 0 0  nmos  L=239.99999143598E-9 W=539.999973625527E-9 
+AD=323.999995669594E-15 AS=194.399997401756E-15 PD=1.74000001607055E-6 
+PS=720.000002729648E-9 M=1 
M266 0 CLK CKON 0  nmos  L=239.99999143598E-9 W=539.999973625527E-9 
+AD=194.399997401756E-15 AS=194.399997401756E-15 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M267 CKON CKO 0 0  nmos  L=239.99999143598E-9 W=539.999973625527E-9 
+AD=194.399997401756E-15 AS=194.399997401756E-15 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M268 0 CKON CKO 0  nmos  L=239.99999143598E-9 W=539.999973625527E-9 
+AD=194.399997401756E-15 AS=194.399997401756E-15 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M269 CKO 1 0 0  nmos  L=239.99999143598E-9 W=539.999973625527E-9 
+AD=194.399997401756E-15 AS=323.999995669594E-15 PD=720.000002729648E-9 
+PS=1.74000001607055E-6 M=1 
   
   
 
.END
