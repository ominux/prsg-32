* # FILE NAME: /HOME/ENGR/LKHWANG/CADENCE/SIMULATION/TOPLEVEL/HSPICES/          
* SCHEMATIC/NETLIST/TOPLEVEL.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON NOV 29 17:17:06 2010
   
* GLOBAL NET DEFINITIONS
.GLOBAL VDD! 
* FILE NAME: PROJECT_TOPLEVEL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TOPLEVEL.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:07 2010.
   
XI23 CLK RESET NET062 NET034 NET061 RESET_G4 
XI16 NET039 NET038 NET33 NET036 CLK NET045 NET062 NET034 NET055 NET061 
+CLOCK_G5 
XI13 NET071 NET066 INV_1 
XI19 NET036 NET046 INV_1 
XI20 NET039 NET0102 INV_1 
XI15 OUT NET026 INV_1 
XI21 NET038 NET082 INV_1 
XI22 NET33 NET087 INV_1 
XI14 NET066 OUT INV_1 
XI12 NET045 NET12 NET071 NET055 TX_GATE_G2 
XI11 NET055 NET16 NET071 NET045 TX_GATE_G2 
XI7 NET11 NET079 NET9 NET12 XOR_G6 
XI6 NET20 NET13 NET091 NET16 XOR_G6 
XLTEMP CLK NET026 NET076 NET023 NET034 D_LATCH_G3 
XL2 NET087 NET11 NET079 NET9 NET33 D_LATCH_G3 
XL4 NET046 NET42 NET086 NET11 NET036 D_LATCH_G3 
XL6 NET0102 NET023 NET043 NET42 NET039 D_LATCH_G3 
XL1 NET0102 NET20 NET091 NET13 NET039 D_LATCH_G3 
XL3 NET082 NET25 NET0101 NET20 NET038 D_LATCH_G3 
XL5 NET087 NET023 NET0106 NET25 NET33 D_LATCH_G3 
   
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:06 2010.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_1 A Y 
M0 Y A 0 0  TSMC25DN  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
   
   
   
* FILE NAME: PROJECT_XOR_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: XOR.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:07 2010.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   NB = NB
*                   Y = Y
.SUBCKT XOR_G6 A B NB Y 
M1 Y A NB 0  TSMC25DN  L=240E-9 W=360E-9 AD=216E-15 AS=216E-15 PD=1.92E-6 
+PS=1.92E-6 M=1 
M0 Y A B VDD!  TSMC25DP  L=240E-9 W=720E-9 AD=432E-15 AS=432E-15 PD=2.64E-6 
+PS=2.64E-6 M=1 
XI0 NB A Y B TX_GATE_G2 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS XOR_G6 
* FILE NAME: PROJECT_CLOCK_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: CLOCK.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:07 2010.
   
* TERMINAL MAPPING: ACT1 = ACT1
*                   ACT2 = ACT2
*                   ACT3 = ACT3
*                   ACT4 = ACT4
*                   CLK = CLK
*                   DIV = DIV
*                   RST = RST
*                   NCLK = NCLK
*                   NDIV = NDIV
*                   NRST = NRST
.SUBCKT CLOCK_G5 ACT1 ACT2 ACT3 ACT4 CLK DIV RST NCLK NDIV NRST 
M1 NDIV NRST VDD! VDD!  TSMC25DP  L=240E-9 W=720E-9 AD=432E-15 AS=432E-15 
+PD=2.64E-6 PS=2.64E-6 M=1 
M0 NET046 RST 0 0  TSMC25DN  L=240E-9 W=360E-9 AD=216E-15 AS=216E-15 
+PD=1.92E-6 PS=1.92E-6 M=1 
XI6 NCLK NDIV ACT4 NAND2_1 
XI4 DIV NCLK ACT2 NAND2_1 
XI5 CLK NDIV ACT3 NAND2_1 
XI3 CLK DIV ACT1 NAND2_1 
XI2 CLK NCLK INV_2 
XI1 CLK NET8 NDIV DIV NCLK D_LATCH_G3 
XI0 NCLK NDIV NET046 NET8 CLK D_LATCH_G3 
   
   
* FILE NAME: NCSU_DIGITAL_PARTS_NAND2_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: NAND2.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:06 2010.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   Y = Y
.SUBCKT NAND2_1 A B Y 
M0 NET9 B 0 0  TSMC25DN  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
M1 Y A NET9 0  TSMC25DN  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
M2 Y A VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
M3 Y B VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS NAND2_1 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:06 2010.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_2 A Y 
M0 Y A 0 0  TSMC25DN  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_2 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS CLOCK_G5 
* FILE NAME: PROJECT_RESET_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: RESET.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:06 2010.
   
* TERMINAL MAPPING: CLK = CLK
*                   IN = IN
*                   RST = RST
*                   NCLK = NCLK
*                   NRST = NRST
.SUBCKT RESET_G4 CLK IN RST NCLK NRST 
XI7 NRST RST INV_1 
XI6 IN NET8 INV_1 
XI5 NET16 IN NRST NAND2_2 
XI4 NET16 CLK NET20 NCLK NDDYNLATCH_G1 
XI3 NET20 NCLK NET8 CLK NDDYNLATCH_G1 
   
   
* FILE NAME: NCSU_DIGITAL_PARTS_NAND2_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: NAND2.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:06 2010.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   Y = Y
.SUBCKT NAND2_2 A B Y 
M0 NET9 B 0 0  TSMC25DN  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
M1 Y A NET9 0  TSMC25DN  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
M2 Y A VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
M3 Y B VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS NAND2_2 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:06 2010.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_1 A Y 
M0 Y A 0 0  TSMC25DN  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS RESET_G4 
* FILE NAME: PROJECT_NDDYNLATCH_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: NDDYNLATCH.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:06 2010.
   
* TERMINAL MAPPING: Q = Q
*                   READ = READ
*                   ND = ND
*                   NREAD = NREAD
.SUBCKT NDDYNLATCH_G1 Q READ ND NREAD 
M3 NET9 ND VDD! VDD!  TSMC25DP  L=240E-9 W=720E-9 AD=432E-15 AS=432E-15 
+PD=2.64E-6 PS=2.64E-6 M=1 
M2 Q NREAD NET9 VDD!  TSMC25DP  L=240E-9 W=720E-9 AD=432E-15 AS=432E-15 
+PD=2.64E-6 PS=2.64E-6 M=1 
M1 Q READ NET16 0  TSMC25DN  L=240E-9 W=360E-9 AD=216E-15 AS=216E-15 
+PD=1.92E-6 PS=1.92E-6 M=1 
M0 NET16 ND 0 0  TSMC25DN  L=240E-9 W=360E-9 AD=216E-15 AS=216E-15 PD=1.92E-6 
+PS=1.92E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS NDDYNLATCH_G1 
* FILE NAME: PROJECT_D_LATCH_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: D_LATCH.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:07 2010.
   
* TERMINAL MAPPING: CLK = CLK
*                   D = D
*                   Q = Q
*                   QB = QB
*                   NCLK = NCLK
.SUBCKT D_LATCH_G3 CLK D Q QB NCLK 
XI3 QB Q INV_1 
XI2 Q QB INV_2 
XI1 CLK D Q NCLK TX_GATE_G2 
   
   
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:06 2010.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_1 A Y 
M0 Y A 0 0  TSMC25DN  L=(600E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC25DP  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:06 2010.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_2 A Y 
M0 Y A 0 0  TSMC25DN  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_2 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS D_LATCH_G3 
* FILE NAME: PROJECT_TX_GATE_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TX_GATE.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV 29 17:17:07 2010.
   
* TERMINAL MAPPING: CLK = CLK
*                   L = L
*                   R = R
*                   NCLK = NCLK
.SUBCKT TX_GATE_G2 CLK L R NCLK 
M1 L CLK R 0  TSMC25DN  L=240E-9 W=360E-9 AD=216E-15 AS=216E-15 PD=1.92E-6 
+PS=1.92E-6 M=1 
M0 L NCLK R VDD!  TSMC25DP  L=240E-9 W=720E-9 AD=432E-15 AS=432E-15 PD=2.64E-6 
+PS=2.64E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TX_GATE_G2 

vVDD VDD! 0 DC 2.5

vCLK CLK 0 pulse(0 2.5 0.5ns 150ps 150ps 350ps 1ns)

vRST Reset 0 pulse(2.5 0 0.5ns 150ps 150ps 23.35ns 24ns)

   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
   
* INCLUDE FILES
   
   
   
* END OF NETLIST
.TEMP    25.0000    
.OP
.save
.option list post=2
.tran 0.01p 24n
.measure tran avgpwr AVG power from=0ns to=100ns
.END
