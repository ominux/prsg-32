* GLOBAL NET DEFINITIONS
.GLOBAL VDD! 
* FILE NAME: PROJECT_TOPLEVEL_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TOPLEVEL.
* GENERATED FOR: HSPICES.
   
XI16 NET039 NET038 NET33 NET036 CLK NET045 NET034 NET055 CLOCK_G3 
XI19 NET039 NET046 INV_1 
XI20 NET038 NET0102 INV_1 
XI15 OUT NET026 INV_1 
XI21 NET33 NET082 INV_1 
XI22 NET036 NET087 INV_1 
XI13 NET071 NET066 INV_1 
XI14 NET066 OUT INV_1 
XI12 NET045 NET12 NET071 NET055 TX_GATE_G1 
XI11 NET055 NET16 NET071 NET045 TX_GATE_G1 
XI7 NET11 NET079 NET9 NET12 XOR_G4 
XI6 NET20 NET13 NET091 NET16 XOR_G4 
XI10 CLK NET026 NET076 NET023 NET034 D_LATCH_G2 
XI5 NET082 NET11 NET079 NET9 NET33 D_LATCH_G2 
XI4 NET087 NET42 NET086 NET11 NET036 D_LATCH_G2 
XI3 NET082 NET023 NET043 NET42 NET33 D_LATCH_G2 
XI2 NET046 NET20 NET091 NET13 NET039 D_LATCH_G2 
XI1 NET0102 NET25 NET0101 NET20 NET038 D_LATCH_G2 
XI0 NET046 NET023 NET0106 NET25 NET039 D_LATCH_G2 
   
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_1 A Y 
M0 Y A 0 0  TSMC25DN  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
   
   
   
* FILE NAME: PROJECT_XOR_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: XOR.
* GENERATED FOR: HSPICES.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   NB = NB
*                   Y = Y
.SUBCKT XOR_G4 A B NB Y 
M1 Y A 0 0  TSMC25DN  L=240E-9 W=360E-9 AD=216E-15 AS=216E-15 PD=1.92E-6 
+PS=1.92E-6 M=1 
M0 Y A VDD! VDD!  TSMC25DP  L=240E-9 W=720E-9 AD=432E-15 AS=432E-15 PD=2.64E-6 
+PS=2.64E-6 M=1 
XI0 NB A Y B TX_GATE_G1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS XOR_G4 
* FILE NAME: PROJECT_CLOCK_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: CLOCK.
* GENERATED FOR: HSPICES.
   
* TERMINAL MAPPING: ACT1 = ACT1
*                   ACT2 = ACT2
*                   ACT3 = ACT3
*                   ACT4 = ACT4
*                   CLK = CLK
*                   DIV = DIV
*                   NCLK = NCLK
*                   NDIV = NDIV
.SUBCKT CLOCK_G3 ACT1 ACT2 ACT3 ACT4 CLK DIV NCLK NDIV 
XI6 NCLK NDIV ACT4 NAND2_1 
XI4 DIV NCLK ACT2 NAND2_1 
XI5 CLK NDIV ACT3 NAND2_1 
XI3 CLK DIV ACT1 NAND2_1 
XI2 CLK NCLK INV_2 
XI1 CLK NET8 NDIV DIV NCLK D_LATCH_G2 
XI0 NCLK NDIV NET046 NET8 CLK D_LATCH_G2 
   
   
* FILE NAME: NCSU_DIGITAL_PARTS_NAND2_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: NAND2.
* GENERATED FOR: HSPICES.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   Y = Y
.SUBCKT NAND2_1 A B Y 
M0 NET9 B 0 0  TSMC25DN  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
M1 Y A NET9 0  TSMC25DN  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
M2 Y A VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
M3 Y B VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS NAND2_1 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_2 A Y 
M0 Y A 0 0  TSMC25DN  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_2 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS CLOCK_G3 
* FILE NAME: PROJECT_D_LATCH_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: D_LATCH.
* GENERATED FOR: HSPICES.
   
* TERMINAL MAPPING: CLK = CLK
*                   D = D
*                   Q = Q
*                   QB = QB
*                   NCLK = NCLK
.SUBCKT D_LATCH_G2 CLK D Q QB NCLK 
XI3 QB Q INV_1 
XI2 Q QB INV_2 
XI1 CLK D Q NCLK TX_GATE_G1 
   
   
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_1 A Y 
M0 Y A 0 0  TSMC25DN  L=(600E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_1 
* FILE NAME: NCSU_DIGITAL_PARTS_INV_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: INV.
* GENERATED FOR: HSPICES.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INV_2 A Y 
M0 Y A 0 0  TSMC25DN  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
M1 Y A VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INV_2 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS D_LATCH_G2 
* FILE NAME: PROJECT_TX_GATE_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: TX_GATE.
* GENERATED FOR: HSPICES.
   
* TERMINAL MAPPING: CLK = CLK
*                   L = L
*                   R = R
*                   NCLK = NCLK
.SUBCKT TX_GATE_G1 CLK L R NCLK 
M1 L CLK R 0  TSMC25DN  L=240E-9 W=360E-9 AD=216E-15 AS=216E-15 PD=1.92E-6 
+PS=1.92E-6 M=1 
M0 L NCLK R VDD!  TSMC25DP  L=240E-9 W=720E-9 AD=432E-15 AS=432E-15 PD=2.64E-6 
+PS=2.64E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS TX_GATE_G1 

vVDD VDD! 0 DC 2.5

vCLK CLK 0 pulse(0 2.5 0.5ns 100ps 100ps 350ps 1ns)


.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
   
* INCLUDE FILES
   
* END OF NETLIST
.TEMP    25.0000    
.OP
.save
.option list post=2
.tran 0.01p 24n
.measure tran avgpwr AVG power from=0ns to=100ns
.END
