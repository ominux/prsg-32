blah

vVDD VDD 0 DC 2.5
vVSS VSS 0 DC 0
vIN IN 0 pulse(2.5 0 1.2ns 100ps 100ps 1.9ns 4ns )

vnCLK nCLK 0 pulse(2.5 0 0.5ns 100ps 100ps 350ps 1ns )
vCLK CLK 0 pulse(0 2.5 0.5ns 100ps 100ps 350ps 1ns )

vnPHI nPHI 0 pulse(0 2.5 .5ns 100ps 100ps 900ps 2ns )
vPHI PHI 0 pulse(2.5 0 .5ns 100ps 100ps 900ps 2ns )

vCON1 P1_1 nPHI DC 0
vCON2 P1_2 CLK DC 0
vCON3 P2_1 nPHI DC 0
vCON4 P2_2 nCLK DC 0
vCON5 P3_1 PHI DC 0
vCON6 P3_2 CLK DC 0
vCON7 P4_1 PHI DC 0
vCON8 P4_2 nCLK DC 0
vCON9 IN D6 DC 0
vCON10 IN D5 DC 0

vnRST nRSTIN 0 pulse(2.5 0 0ns 100ps 100ps 0.4ns 80ns )
vRST RSTIN 0 pulse(0 2.5 0ns 100ps 100ps 0.4ns 80ns)

* Reset transistors for latches.

M103 Q1 nRSTIN VDD VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 

M104 Q6 nRSTIN VDD VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 

M105 nQ3 RSTIN VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1

M106 nQ4 RSTIN VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1

*end of reset transistors


.OPTION list post=2   
.tran 0.01p 24n
.measure tran avgpwr AVG power from=0ns to=100ns
   
M43 VDD 8 6 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=475.200011718774E-15 PD=1.91999993148784E-6 
+PS=2.04000002668181E-6 M=1 
M44 VDD 7 5 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=475.200011718774E-15 PD=1.91999993148784E-6 
+PS=2.04000002668181E-6 M=1 
M45 4 2 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=475.200011718774E-15 AS=432.000003261143E-15 PD=2.04000002668181E-6 
+PS=1.91999993148784E-6 M=1 
M46 3 1 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=475.200011718774E-15 AS=432.000003261143E-15 PD=2.04000002668181E-6 
+PS=1.91999993148784E-6 M=1 
M47 Q2 8 42 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M48 42 NQ4 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M49 NQ4 7 41 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M50 41 Q6 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M51 Q6 1 40 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M52 40 D6 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M53 VDD D5 39 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M54 39 8 Q5 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M55 VDD Q5 38 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M56 38 2 NQ3 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M57 VDD NQ3 37 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M58 37 1 Q1 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M59 7 P2_2 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=388.799994803513E-15 PD=2.27999998969608E-6 
+PS=720.000002729648E-9 M=1 
M60 8 P1_2 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=388.799994803513E-15 PD=2.27999998969608E-6 
+PS=720.000002729648E-9 M=1 
M61 VDD P1_1 8 VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M62 VDD P2_1 7 VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M63 2 P4_2 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=388.799994803513E-15 PD=2.27999998969608E-6 
+PS=720.000002729648E-9 M=1 
M64 1 P3_2 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=388.799994803513E-15 PD=2.27999998969608E-6 
+PS=720.000002729648E-9 M=1 
M65 VDD P3_1 1 VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M66 VDD P4_1 2 VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M67 Q2 6 16 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M68 16 NQ4 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M69 NQ4 5 15 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M70 15 Q6 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M71 Q6 3 14 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M72 14 D6 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M73 VSS D5 13 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M74 13 6 Q5 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M75 VSS Q5 12 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M76 12 4 NQ3 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M77 VSS NQ3 11 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M78 11 3 Q1 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M79 VSS P1_2 18 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=129.599998267838E-15 PD=1.7999999499807E-6 
+PS=720.000002729648E-9 M=1 
M80 VSS P2_2 17 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=129.599998267838E-15 PD=1.7999999499807E-6 
+PS=720.000002729648E-9 M=1 
M81 18 P1_1 8 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=129.599998267838E-15 AS=273.599990319867E-15 PD=720.000002729648E-9 
+PS=1.7999999499807E-6 M=1 
M82 17 P2_1 7 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=129.599998267838E-15 AS=273.599990319867E-15 PD=720.000002729648E-9 
+PS=1.7999999499807E-6 M=1 
M83 VSS 8 6 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M84 VSS 7 5 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M85 4 2 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M86 3 1 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M87 1 P3_2 9 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=129.599998267838E-15 PD=1.7999999499807E-6 
+PS=720.000002729648E-9 M=1 
M88 2 P4_2 10 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=129.599998267838E-15 PD=1.7999999499807E-6 
+PS=720.000002729648E-9 M=1 
M89 10 P4_1 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=129.599998267838E-15 AS=273.599990319867E-15 PD=720.000002729648E-9 
+PS=1.7999999499807E-6 M=1 
M90 9 P3_1 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=129.599998267838E-15 AS=273.599990319867E-15 PD=720.000002729648E-9 
+PS=1.7999999499807E-6 M=1 
   
   
   
   
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
   
* INCLUDE FILES
   
   
.END
