

***********LATCHES****************

*Using Static Latches
*X1 nQ3 Q1 READP3 nREADP3 VDD 0 nDLATCH
*X3 Q5 nQ3 READP4 nREADP4 VDD 0 nDLATCH
*X5 nQT Q5 READP1 nREADP1 VDD 0 nDLATCH
*X2 nQ4 Q2 READP1 nREADP1 VDD 0 nDLATCH
*X4 Q6 nQ4 READP2 nREADP2 VDD 0 nDLATCH
*X6 nQT Q6 READP3 nREADP3 VDD 0 nDLATCH
*XT IN nQT nCLK CLK VDD 0 nDLATCH

*Using Dynamic Latches
X1 nQ3 Q1 READP3 nREADP3 VDD 0 nDDYNLATCH
X3 Q5 nQ3 READP4 nREADP4 VDD 0 nDDYNLATCH
X5 nQT Q5 READP1 nREADP1 VDD 0 nDDYNLATCH
X2 nQ4 Q2 READP1 nREADP1 VDD 0 nDDYNLATCH
X4 Q6 nQ4 READP2 nREADP2 VDD 0 nDDYNLATCH
X6 nQT Q6 READP3 nREADP3 VDD 0 nDDYNLATCH
XT IN nQT nCLK CLK VDD 0 nDDYNLATCH

XRST RSTIN CLK nCLK RST nRST VDD 0 RESET

**************LATCH CLOCKING***************

X3c CLK nPHI nREADP3 READP3 VDD 0 NAND2_CLK
X4c nCLK nPHI nREADP4 READP4 VDD 0 NAND2_CLK
X1c CLK PHI nREADP1 READP1 VDD 0 NAND2_CLK
X2c nCLK PHI nREADP2 READP2 VDD 0 NAND2_CLK

.subckt nDLATCH nD Q READ nREAD VDD VSS

MTP1 nD nREAD QB VDD TSMC25DP L=240E-9 W=720E-9 
+AD=432E-15 AS=432E-15 PD=1.92E-6 
+PS=1.92E-6 M=1
MTN1 nD READ QB VSS TSMC25DN L=240E-9 W=360E-9 
+AD=216E-15 AS=216E-15 PD=1.56E-6 
+PS=1.56E-6 M=1 

MPI1 Q QB VDD VDD TSMC25DP L=240E-9 W=720E-9 
+AD=432E-15 AS=432E-15 PD=1.92E-6 
+PS=1.92E-6 M=1
MNI1 Q QB VSS VSS TSMC25DN L=240E-9 W=360E-9 
+AD=216E-15 AS=216E-15 PD=1.56E-6 
+PS=1.56E-6 M=1

MPI2 QB Q VDD VDD TSMC25DP L=240E-9 W=360E-9 
+AD=432E-15 AS=432E-15 PD=1.92E-6 
+PS=1.92E-6 M=1 
MNI2 QB Q VSS VSS TSMC25DN L=600E-9 W=360E-9 
+AD=216E-15 AS=216E-15 PD=1.56E-6 
+PS=1.56E-6 M=1
.ends

.subckt nDDYNLATCH nD Q READ nREAD VDD VSS

MPgate Q nREAD INTP VDD TSMC25DP L=240E-9 W=720E-9 
+AD=432E-15 AS=432E-15 PD=1.92E-6 
+PS=1.92E-6 M=1
MNgate Q READ INTN VSS TSMC25DN L=240E-9 W=360E-9 
+AD=216E-15 AS=216E-15 PD=1.56E-6 
+PS=1.56E-6 M=1

MPdata INTP nD VDD VDD TSMC25DP L=240E-9 W=720E-9 
+AD=432E-15 AS=432E-15 PD=1.92E-6 
+PS=1.92E-6 M=1
MNdata INTN nD VSS VSS TSMC25DN L=240E-9 W=360E-9 
+AD=216E-15 AS=216E-15 PD=1.56E-6 
+PS=1.56E-6 M=1

.ends

.subckt NAND2_CLK A B OUT nOUT VDD VSS

MPnand1 OUT A VDD VDD TSMC25DP L=240E-9 W=1.08E-6 
+AD=648E-15 AS=648E-15 PD=2.28E-6 
+PS=2.28E-6 M=1
MPnand2 OUT B VDD VDD TSMC25DP L=240E-9 W=1.08E-6 
+AD=648E-15 AS=648E-15 PD=2.28E-6 
+PS=2.28E-6 M=1

MNnand1 OUT A 1 VSS TSMC25DN L=240E-9 W=360E-9 
+AD=216E-15 AS=216E-15 PD=1.56E-6 
+PS=1.56E-6 M=1
MNnand2 1 B VSS VSS TSMC25DN L=240E-9 W=360E-9 
+AD=216E-15 AS=216E-15 PD=1.56E-6 
+PS=1.56E-6 M=1

MNI nOUT OUT VSS VSS TSMC25DN L=240E-9 W=360E-9 
+AD=216E-15 AS=216E-15 PD=1.56E-6 
+PS=1.56E-6 M=1
MPI nOUT OUT VDD VDD TSMC25DP L=240E-9 W=1.08E-6 
+AD=648E-15 AS=648E-15 PD=2.28E-6 
+PS=2.28E-6 M=1

.ends

.subckt RESET IN CLK nCLK RST nRST VDD VSS

MPI1 nIN IN VDD VDD TSMC25DP L=240E-9 W=720E-9 
+AD=432E-15 AS=432E-15 PD=1.92E-6 
+PS=1.92E-6 M=1
MNI1 nIN IN VSS VSS TSMC25DN L=240E-9 W=360E-9 
+AD=216E-15 AS=216E-15 PD=1.56E-6 
+PS=1.56E-6 M=1

MPI2 RST nRST VDD VDD TSMC25DP L=240E-9 W=720E-9 
+AD=432E-15 AS=432E-15 PD=1.92E-6 
+PS=1.92E-6 M=1
MNI2 RST nRST VSS VSS TSMC25DN L=240E-9 W=360E-9 
+AD=216E-15 AS=216E-15 PD=1.56E-6 
+PS=1.56E-6 M=1

MPnand1 nRST Qr VDD VDD TSMC25DP L=240E-9 W=720E-9 
+AD=432E-15 AS=432E-15 PD=1.92E-6 
+PS=1.92E-6 M=1
MPnand2 nRST IN VDD VDD TSMC25DP L=240E-9 W=720E-9 
+AD=432E-15 AS=432E-15 PD=1.92E-6 
+PS=1.92E-6 M=1

MNnand1 nRST Qr 1 VSS TSMC25DN L=240E-9 W=720E-9 
+AD=432E-15 AS=432E-15 PD=1.92E-6 
+PS=1.92E-6 M=1
MNnand2 1 IN VSS VSS TSMC25DN L=240E-9 W=720E-9 
+AD=432E-15 AS=432E-15 PD=1.92E-6 
+PS=1.92E-6 M=1

Xf nIN Qf nCLK CLK VDD 0 nDDYNLATCH
Xr Qf Qr  CLK nCLK VDD 0 nDDYNLATCH

.ends

.subckt CKDIV CK2 nCK2 CLK nCLK VDD VSS 

x1 nCK2 Q NCLK CLK VDD VSS nDLATCH
x2 Q CK2 CLK nCLK VDD VSS nDLATCH

MTP1 nCK2 CK2 VDD VDD TSMC25DP L=240E-9 W=720E-9 
+AD=432E-15 AS=432E-15 PD=1.92E-6 
+PS=1.92E-6 M=1
MTN1 nCK2 CK2 VSS VSS TSMC25DN L=240E-9 W=360E-9 
+AD=216E-15 AS=216E-15 PD=1.56E-6 
+PS=1.56E-6 M=1 

.ends

vVDD VDD 0 DC 2.5
vIN IN 0 pulse(2.5 0 1ns 100ps 100ps 1.9ns 4ns )

vnCLK nCLK 0 pulse(2.5 0 0.5ns 100ps 100ps 350ps 1ns )
vCLK CLK 0 pulse(0 2.5 0.5ns 100ps 100ps 350ps 1ns )

vnPHI nPHI 0 pulse(0 2.5 .5ns 100ps 100ps 900ps 2ns )
vPHI PHI 0 pulse(2.5 0 .5ns 100ps 100ps 900ps 2ns )

vRST RSTIN 0 pulse(2.5 0 1ns 100ps 100ps 3ns 8ns )

.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 

.OPTION list post=2   
.tran 0.01p 24n
.measure tran avgpwr AVG power from=0ns to=100ns

.END

