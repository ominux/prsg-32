blah

vVDD VDD 0 DC 2.5
vVSS VSS 0 DC 0
vIN IN 0 pulse(2.5 0 1.2ns 100ps 100ps 1.9ns 4ns )

*vnCLK nCLK 0 pulse(2.5 0 0.6ns 100ps 100ps .4ns 1ns )
vCLK CLK 0 pulse(0 2.5 0.5ns 100ps 100ps 0.4ns 1ns )

*vnPHI nPHI 0 pulse(0 2.5 .5ns 100ps 100ps 900ps 2ns )
*vPHI PHI 0 pulse(2.5 0 .5ns 100ps 100ps 900ps 2ns )

.OPTION list post=2   
.tran 0.01p 100n
.measure tran avgpwr AVG power from=0ns to=100ns

MPI1 CKO CLK VDD VDD pmos  L=239.99999143598E-9 W=1.0800000054593E-6 
+AD=648.000006522286E-15 AS=648.000006522286E-15 PD=2.28000004790432E-6 
+PS=2.28000004790432E-6 M=1   
MNI1 CKO CLK 0 0 nmos  L=239.99999143598E-9 W=540.000002729648E-9 
+AD=324.199996535675E-15 AS=324.199996535675E-15 PD=1740.000002729648E-9 
+PS=1740.000002729648E-9 M=1 
MPI2 1 CLK VDD VDD pmos L=239.99999143598E-9 W=1.0800000054593E-6 
+AD=648.000006522286E-15 AS=648.000006522286E-15 PD=2.28000004790432E-6 
+PS=2.28000004790432E-6 M=1 
MNI2 1 CLK 0 0 nmos  L=239.99999143598E-9 W=540.000002729648E-9 
+AD=324.199996535675E-15 AS=324.199996535675E-15 PD=1740.000002729648E-9 
+PS=1740.000002729648E-9 M=1  
MPI3 nCKO 1 VDD VDD pmos  L=239.99999143598E-9 W=1.0800000054593E-6 
+AD=648.000006522286E-15 AS=648.000006522286E-15 PD=2.28000004790432E-6 
+PS=2.28000004790432E-6 M=1     
MNI3 nCKO 1 0 0 nmos  L=239.99999143598E-9 W=540.000002729648E-9 
+AD=324.199996535675E-15 AS=324.199996535675E-15 PD=1740.000002729648E-9 
+PS=1740.000002729648E-9 M=1   
MPI4 nCKO CKO VDD VDD pmos  L=239.99999143598E-9 W=1.0800000054593E-6 
+AD=648.000006522286E-15 AS=648.000006522286E-15 PD=2.28000004790432E-6 
+PS=2.28000004790432E-6 M=1  
MNI4 nCKO CKO 0 0 nmos  L=239.99999143598E-9 W=540.000002729648E-9 
+AD=324.199996535675E-15 AS=324.199996535675E-15 PD=1740.000002729648E-9 
+PS=1740.000002729648E-9 M=1 
MPI5 CKO nCKO VDD VDD pmos  L=239.99999143598E-9 W=1.0800000054593E-6 
+AD=648.000006522286E-15 AS=648.000006522286E-15 PD=2.28000004790432E-6 
+PS=2.28000004790432E-6 M=1 
MNI5 CKO nCKO 0 0 nmos L=239.99999143598E-9 W=540.000002729648E-9 
+AD=324.199996535675E-15 AS=324.199996535675E-15 PD=1740.000002729648E-9 
+PS=1740.000002729648E-9 M=1 



x1  CKO OUT4 OUT3 OUT1 VDD VSS NAND3
x2  nCKO  OUT1 OUT4 OUT2 VDD VSS NAND3
x3  CKO  OUT2 OUT1 OUT3 VDD VSS NAND3
x4  nCKO  OUT3 OUT2 OUT4 VDD VSS NAND3
 



.subckt NAND3 A B C OUT VDD VSS
M45 OUT A VDD VDD  pmos  L=239.99999143598E-9 W=2.88000001091859E-6 
+AD=1.72800001304457E-12 AS=1.72800001304457E-12 PD=4.08000005336362E-6 
+PS=4.08000005336362E-6 M=1 
*M46 OUT B VDD VDD  pmos  L=239.99999143598E-9 W=2.16000001091859E-6 
*+AD=1.72800001304457E-12 AS=1.72800001304457E-12 PD=4.08000005336362E-6 
*+PS=4.08000005336362E-6 M=1 
*M47 OUT C VDD VDD  pmossvn   L=239.99999143598E-9 W=1.8000000054593E-6 
*+AD=1080.000006522286E-15 AS=1080.000006522286E-15 PD=3.00000004790432E-6 
*+PS=2.64000004790432E-6 M=1 

M48 1 A VSS VSS  nmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M49 1 B 2 VSS  nmos  L=239.99999143598E-9 W=1.07999994725105E-6 +AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M50 OUT C 2 VSS  nmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
.ends
   
*.lib "$CDK_DIR/models/hspice/public/publicModel/nmos" NMOS 
*.lib "$CDK_DIR/models/hspice/public/publicModel/pmos" PMOS 


.lib 'models25.txt' SS
* INCLUDE FILES
   
   
.END

vcon0A nCLK 0 DC 0
vCON1 P1_1 nPHI DC 0
vCON2 P1_2 CLK DC 0
vCON3 P2_1 nPHI DC 0
vCON4 P2_2 nCLK DC 0
vCON5 P3_1 PHI DC 0
vCON6 P3_2 CLK DC 0
vCON7 P4_1 PHI DC 0
vCON8 P4_2 nCLK DC 0
vCON9 IN D6 DC 0
vCON10 IN D5 DC 0

vnRST nRSTIN 0 pulse(2.5 0 0ns 100ps 100ps 0.4ns 80ns )
vRST RSTIN 0 pulse(0 2.5 0ns 100ps 100ps 0.4ns 80ns)

* Clock division circuit (should be swapped?)
XPHI CLK nclk nPHI pu vdd clk_div
XnPHI CLK nclk PHI pd vdd clk_div

M101 pd RSTIN VSS VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1

M102 pu nRSTIN VDD VDD  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 

* Reset transistors for latches.


M103 Q1 nRSTIN VDD VDD  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 

M104 Q6 nRSTIN VDD VDD  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 

M105 nQ3 RSTIN VSS VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1

M106 nQ4 RSTIN VSS VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1




.OPTION list post=2   
.tran 0.01p 24n
.measure tran avgpwr AVG power from=0ns to=100ns
   
M43 VDD 8 6 VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=475.200011718774E-15 PD=1.91999993148784E-6 
+PS=2.04000002668181E-6 M=1 
M44 VDD 7 5 VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=475.200011718774E-15 PD=1.91999993148784E-6 
+PS=2.04000002668181E-6 M=1 
M45 4 2 VDD VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=475.200011718774E-15 AS=432.000003261143E-15 PD=2.04000002668181E-6 
+PS=1.91999993148784E-6 M=1 
M46 3 1 VDD VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=475.200011718774E-15 AS=432.000003261143E-15 PD=2.04000002668181E-6 
+PS=1.91999993148784E-6 M=1 
M47 Q2 8 42 VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M48 42 NQ4 VDD VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M49 NQ4 7 41 VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M50 41 Q6 VDD VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M51 Q6 1 40 VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M52 40 D6 VDD VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M53 VDD D5 39 VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M54 39 8 Q5 VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M55 VDD Q5 38 VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M56 38 2 NQ3 VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M57 VDD NQ3 37 VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M58 37 1 Q1 VDD  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M59 7 P2_2 VDD VDD  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=388.799994803513E-15 PD=2.27999998969608E-6 
+PS=720.000002729648E-9 M=1 
M60 8 P1_2 VDD VDD  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=388.799994803513E-15 PD=2.27999998969608E-6 
+PS=720.000002729648E-9 M=1 
M61 VDD P1_1 8 VDD  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M62 VDD P2_1 7 VDD  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M63 2 P4_2 VDD VDD  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=388.799994803513E-15 PD=2.27999998969608E-6 
+PS=720.000002729648E-9 M=1 
M64 1 P3_2 VDD VDD  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=388.799994803513E-15 PD=2.27999998969608E-6 
+PS=720.000002729648E-9 M=1 
M65 VDD P3_1 1 VDD  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M66 VDD P4_1 2 VDD  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M67 Q2 6 16 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M68 16 NQ4 VSS VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M69 NQ4 5 15 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M70 15 Q6 VSS VSS o nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M71 Q6 3 14 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M72 14 D6 VSS VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M73 VSS D5 13 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M74 13 6 Q5 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M75 VSS Q5 12 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M76 12 4 NQ3 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M77 VSS NQ3 11 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M78 11 3 Q1 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M79 VSS P1_2 18 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=129.599998267838E-15 PD=1.7999999499807E-6 
+PS=720.000002729648E-9 M=1 
M80 VSS P2_2 17 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=129.599998267838E-15 PD=1.7999999499807E-6 
+PS=720.000002729648E-9 M=1 
M81 18 P1_1 8 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=129.599998267838E-15 AS=273.599990319867E-15 PD=720.000002729648E-9 
+PS=1.7999999499807E-6 M=1 
M82 17 P2_1 7 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=129.599998267838E-15 AS=273.599990319867E-15 PD=720.000002729648E-9 
+PS=1.7999999499807E-6 M=1 
M83 VSS 8 6 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.799999949980o7E-6 M=1 
M84 VSS 7 5 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M85 4 2 VSS VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M86 3 1 VSS VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M87 1 P3_2 9 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=129.599998267838E-15 PD=1.7999999499807E-6 
+PS=720.000002729648E-9 M=1 
M88 2 P4_2 10 VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=129.599998267838E-15 PD=1.7999999499807E-6 
+PS=720.000002729648E-9 M=1 
M89 10 P4_1 VSS VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=129.599998267838E-15 AS=273.599990319867E-15 PD=720.000002729648E-9 
+PS=1.7999999499807E-6 M=1 
M90 9 P3_1 VSS VSS  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=129.599998267838E-15 AS=273.599990319867E-15 PD=720.000002729648E-9 
+PS=1.7999999499807E-6 M=1   
   
   
  
.subckt clk_div clk nclk DIVCLK set vdd
C6 0 1  30.7296E-18 M=1.0 
C7 SET 0  42.6024E-18 M=1.0 
C8 VDD 1  44.6976E-18 M=1.0 
C9 VDD SET  30.0312E-18 M=1.0 
C10 DIVCLK 0  37.7136E-18 M=1.0 
C11 DIVCLK VDD  34.92E-18 M=1.0 
C12 CLK 0  41.904E-18 M=1.0 
C13 CLK VDD  32.1264E-18 M=1.0 
C14 NCLK 0  40.5072E-18 M=1.0 
C15 NCLK VDD  36.3168E-18 M=1.0 
C16 0 1  51.2496E-18 M=1.0 
C17 SET 0  78.7896E-18 M=1.0 
C18 VDD 1  71.616E-18 M=1.0 
C19 VDD 0  335.2512E-18 M=1.0 
C20 VDD SET  78.8376E-18 M=1.0 
C21 DIVCLK 0  89.2704E-18 M=1.0 
C22 DIVCLK VDD  63.9312E-18 M=1.0 
C23 CLK 0  77.208E-18 M=1.0 
C24 NCLK 5  25.92E-18 M=1.0 
C25 NCLK 0  86.2848E-18 M=1.0 
C26 NCLK VDD  106.6152E-18 M=1.0 
C27 DIVCLK 1  100.5336E-18 M=1.0 
C28 DIVCLK SET  100.5408E-18 M=1.0 
C29 DIVCLK VDD  367.524E-18 M=1.0 
C30 CLK 0  1.194744E-15 M=1.0 
C31 CLK VDD  475.6848E-18 M=1.0 
C32 CLK DIVCLK  36.864E-18 M=1.0 
C33 NCLK 1  122.184E-18 M=1.0 
C34 NCLK 0  283.6728E-18 M=1.0 
C35 NCLK DIVCLK  90.648E-18 M=1.0 
M36 1 CLK 4 VDD  pmos  L=239.99999143598E-9 W=2.88000001091859E-6 
+AD=1.72800001304457E-12 AS=1.72800001304457E-12 PD=4.08000005336362E-6 
+PS=4.08000005336362E-6 M=1  
M37 4 DIVCLK VDD VDD  pmos  L=239.99999143598E-9 W=2.88000001091859E-6 
+AD=1.72800001304457E-12 AS=1.72800001304457E-12 PD=4.08000005336362E-6 
+PS=4.08000005336362E-6 M=1  
M38 SET NCLK 5 VDD  pmos  L=239.99999143598E-9 W=2.88000001091859E-6 
+AD=1.72800001304457E-12 AS=1.72800001304457E-12 PD=4.08000005336362E-6 
+PS=4.08000005336362E-6 M=1 
M39 5 1 VDD VDD  pmos  L=239.99999143598E-9 W=2.88000001091859E-6 
+AD=1.72800001304457E-12 AS=1.72800001304457E-12 PD=4.08000005336362E-6 
+PS=4.08000005336362E-6 M=1 
M40 DIVCLK SET VDD VDD  pmos  L=239.99999143598E-9 W=2.88000001091859E-6 
+AD=1.72800001304457E-12 AS=1.72800001304457E-12 PD=4.08000005336362E-6 
+PS=4.08000005336362E-6 M=1 
M41 1 NCLK 2 0  nmos  L=239.99999143598E-9 W=1.4400000054593E-6 
+AD=864.000006522286E-15 AS=864.000006522286E-15 PD=2.64000004790432E-6 
+PS=2.64000004790432E-6 M=1  
M42 2 DIVCLK 0 0  nmos  L=239.99999143598E-9 W=1.4400000054593E-6 
+AD=864.000006522286E-15 AS=864.000006522286E-15 PD=2.64000004790432E-6 
+PS=2.64000004790432E-6 M=1  
M43 SET CLK 3 0  nmos  L=239.99999143598E-9 W=1.4400000054593E-6 
+AD=864.000006522286E-15 AS=864.000006522286E-15 PD=2.64000004790432E-6 
+PS=2.64000004790432E-6 M=1  
M44 3 1 0 0  nmos  L=239.99999143598E-9 W=1.4400000054593E-6 
+AD=864.000006522286E-15 AS=864.000006522286E-15 PD=2.64000004790432E-6 
+PS=2.64000004790432E-6 M=1 
M45 DIVCLK SET 0 0  nmos  L=239.99999143598E-9 W=1.4400000054593E-6 
+AD=864.000006522286E-15 AS=864.000006522286E-15 PD=2.64000004790432E-6 
+PS=2.64000004790432E-6 M=1 
.ends
