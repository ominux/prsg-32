blah

vVDD VDD 0 DC 2.5
vVSS VSS 0 DC 0
vIN IN 0 pulse(2.5 0 1.2ns 100ps 100ps 1.9ns 4ns )

*vnCLK nCLK 0 pulse(2.5 0 0.5ns 100ps 100ps 350ps 1ns )
vCK CK 0 pulse(0 2.5 0.5ns 100ps 100ps 350ps 1ns )

*vnPHI nPHI 0 pulse(0 2.5 .5ns 100ps 100ps 900ps 2ns )
*vPHI PHI 0 pulse(2.5 0 .5ns 100ps 100ps 900ps 2ns )

vCON1 P11 nPHI DC 0
vCON2 P12 CLK DC 0
vCON3 P21 nPHI DC 0
vCON4 P22 nCLK DC 0
vCON5 P31 PHI DC 0
vCON6 P32 CLK DC 0
vCON7 P41 PHI DC 0
vCON8 P42 nCLK DC 0
vCON9 IN D6 DC 0
vCON10 IN D5 DC 0

vRST RSTIN 0 pulse(2.5 0 1ns 100ps 100ps 3ns 8ns )

.OPTION list post=2   
.tran 0.01p 24n
.measure tran avgpwr AVG power from=0ns to=100ns

x1 CK CLK NCLK PHI VDD! 0 ckmaker
x2 CK CLK NCLK nPHI VDD! 0 ckmaker
x3 CK CLK NCLK PHI VDD! 0 ckmaker
x4 CK CLK NCLK nPHI VDD! 0 ckmaker
   
M43 VDD 8 6 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=475.200011718774E-15 PD=1.91999993148784E-6 
+PS=2.04000002668181E-6 M=1 
M44 VDD 7 5 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=475.200011718774E-15 PD=1.91999993148784E-6 
+PS=2.04000002668181E-6 M=1 
M45 4 2 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=475.200011718774E-15 AS=432.000003261143E-15 PD=2.04000002668181E-6 
+PS=1.91999993148784E-6 M=1 
M46 3 1 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=475.200011718774E-15 AS=432.000003261143E-15 PD=2.04000002668181E-6 
+PS=1.91999993148784E-6 M=1 
M47 NQ4 8 41 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M48 41 Q6 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M49 Q6 7 40 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M50 40 D6 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M51 Q2 2 42 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M52 42 NQ4 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M53 VDD D5 39 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M54 39 2 Q5 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M55 VDD Q5 38 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M56 38 1 NQ3 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M57 VDD NQ3 37 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M58 37 7 Q1 VDD  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M59 8 P22 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=388.799994803513E-15 PD=2.27999998969608E-6 
+PS=720.000002729648E-9 M=1 
M60 7 P31 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=388.799994803513E-15 PD=2.27999998969608E-6 
+PS=720.000002729648E-9 M=1 
M61 VDD P21 8 VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M62 VDD P32 7 VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M63 1 P41 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=388.799994803513E-15 PD=2.27999998969608E-6 
+PS=720.000002729648E-9 M=1 
M64 2 P12 VDD VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=388.799994803513E-15 PD=2.27999998969608E-6 
+PS=720.000002729648E-9 M=1 
M65 VDD P11 2 VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M66 VDD P42 1 VDD  TSMC25DP  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=388.799994803513E-15 AS=647.999991339188E-15 PD=720.000002729648E-9 
+PS=2.27999998969608E-6 M=1 
M67 Q2 4 16 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M68 16 NQ4 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M69 NQ4 6 15 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M70 15 Q6 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M71 Q6 5 14 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M72 14 D6 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M73 VSS D5 13 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M74 13 4 Q5 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M75 VSS Q5 12 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M76 12 3 NQ3 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M77 VSS NQ3 11 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M78 11 5 Q1 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M79 VSS P22 18 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=129.599998267838E-15 PD=1.7999999499807E-6 
+PS=720.000002729648E-9 M=1 
M80 VSS P31 17 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=129.599998267838E-15 PD=1.7999999499807E-6 
+PS=720.000002729648E-9 M=1 
M81 18 P21 8 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=129.599998267838E-15 AS=273.599990319867E-15 PD=720.000002729648E-9 
+PS=1.7999999499807E-6 M=1 
M82 17 P32 7 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=129.599998267838E-15 AS=273.599990319867E-15 PD=720.000002729648E-9 
+PS=1.7999999499807E-6 M=1 
M83 VSS 8 6 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M84 VSS 7 5 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M85 3 1 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M86 4 2 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M87 2 P12 10 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=129.599998267838E-15 PD=1.7999999499807E-6 
+PS=720.000002729648E-9 M=1 
M88 1 P41 9 VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=129.599998267838E-15 PD=1.7999999499807E-6 
+PS=720.000002729648E-9 M=1 
M89 10 P11 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=129.599998267838E-15 AS=273.599990319867E-15 PD=720.000002729648E-9 
+PS=1.7999999499807E-6 M=1 
M90 9 P42 VSS VSS  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=129.599998267838E-15 AS=273.599990319867E-15 PD=720.000002729648E-9 
+PS=1.7999999499807E-6 M=1 

.subckt ckmaker IN CK NCK CKDIV VDD! 0
   
C14 0 3  42.6024E-18 M=1.0 
C15 0 2  30.7296E-18 M=1.0 
C16 0 1  26.19E-18 M=1.0 
C17 VDD! 3  30.0312E-18 M=1.0 
C18 VDD! 2  44.6976E-18 M=1.0 
C19 VDD! 1  40.8564E-18 M=1.0 
C20 CKDIV 0  37.7136E-18 M=1.0 
C21 CKDIV VDD!  34.92E-18 M=1.0 
C22 CK 0  50.2848E-18 M=1.0 
C23 CK VDD!  23.7456E-18 M=1.0 
C24 IN 0  110.3472E-18 M=1.0 
C25 IN VDD!  128.5056E-18 M=1.0 
C26 NCK 0  67.0464E-18 M=1.0 
C27 NCK VDD!  79.6176E-18 M=1.0 
C28 0 3  78.7896E-18 M=1.0 
C29 0 2  51.2496E-18 M=1.0 
C30 0 1  83.9232E-18 M=1.0 
C31 VDD! 3  78.8376E-18 M=1.0 
C32 VDD! 2  71.616E-18 M=1.0 
C33 VDD! 1  94.9392E-18 M=1.0 
C34 VDD! 0  620.3952E-18 M=1.0 
C35 CKDIV 0  89.2704E-18 M=1.0 
C36 CKDIV VDD!  63.9312E-18 M=1.0 
C37 CK 0  156.7344E-18 M=1.0 
C38 CK VDD!  51.2496E-18 M=1.0 
C39 IN 0  99.264E-18 M=1.0 
C40 NCK 13  25.92E-18 M=1.0 
C41 NCK 0  181.6464E-18 M=1.0 
C42 NCK VDD!  254.9568E-18 M=1.0 
C43 NCK 0  719.0952E-18 M=1.0 
C44 NCK VDD!  69.6312E-18 M=1.0 
C45 0 1  258.9168E-18 M=1.0 
C46 VDD! 1  262.4736E-18 M=1.0 
C47 CKDIV 3  100.5408E-18 M=1.0 
C48 CKDIV 2  100.5336E-18 M=1.0 
C49 CKDIV VDD!  367.524E-18 M=1.0 
C50 CK 1  90.648E-18 M=1.0 
C51 IN 1  73.728E-18 M=1.0 
C52 IN 0  2.0609472E-15 M=1.0 
C53 IN VDD!  969.9624E-18 M=1.0 
C54 IN CKDIV  36.864E-18 M=1.0 
C55 NCK 2  122.184E-18 M=1.0 
C56 NCK 1  129.9528E-18 M=1.0 
C57 NCK 0  283.6728E-18 M=1.0 
C58 NCK CKDIV  90.648E-18 M=1.0 
C59 NCK IN  75.4848E-18 M=1.0 
C60 0 1  94.0464E-18 M=1.0 
C61 VDD! 1  79.956E-18 M=1.0 
C62 CK 0  94.1904E-18 M=1.0 
C63 CK VDD!  80.4096E-18 M=1.0 
C64 IN 0  92.3616E-18 M=1.0 
C65 IN VDD!  92.3616E-18 M=1.0 
C66 NCK 0  120.3168E-18 M=1.0 
C67 NCK VDD!  119.37E-18 M=1.0 
M68 VDD! NCK CK VDD!  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=259.199996535675E-15 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M69 CK 1 VDD! VDD!  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=432.000003261143E-15 PD=720.000002729648E-9 
+PS=1.91999993148784E-6 M=1 
M70 1 IN VDD! VDD!  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=259.199996535675E-15 PD=1.91999993148784E-6 
+PS=720.000002729648E-9 M=1 
M71 VDD! IN NCK VDD!  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=259.199996535675E-15 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M72 NCK CK VDD! VDD!  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=259.199996535675E-15 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M73 2 IN 6 VDD!  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M74 6 CKDIV VDD! VDD!  TSMC25DP  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M75 3 NCK 13 VDD!  TSMC25DP  L=239.99999143598E-9 W=1.4400000054593E-6 
+AD=864.000006522286E-15 AS=345.600013450936E-15 PD=2.64000004790432E-6 
+PS=479.999982871959E-9 M=1 
M76 13 2 VDD! VDD!  TSMC25DP  L=239.99999143598E-9 W=1.4400000054593E-6 
+AD=345.600013450936E-15 AS=864.000006522286E-15 PD=479.999982871959E-9 
+PS=2.64000004790432E-6 M=1 
M77 CKDIV 3 VDD! VDD!  TSMC25DP  L=239.99999143598E-9 W=2.88000001091859E-6 
+AD=1.72800001304457E-12 AS=1.72800001304457E-12 PD=4.08000005336362E-6 
+PS=4.08000005336362E-6 M=1 
M78 CK 1 0 0  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=273.599990319867E-15 PD=839.999984236783E-9 
+PS=1.7999999499807E-6 M=1 
M79 1 IN 0 0  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=158.399999388749E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M80 0 IN NCK 0  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=158.399999388749E-15 PD=839.999984236783E-9 
+PS=839.999984236783E-9 M=1 
M81 NCK CK 0 0  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=158.399999388749E-15 PD=839.999984236783E-9 
+PS=839.999984236783E-9 M=1 
M82 0 NCK CK 0  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=158.399999388749E-15 PD=839.999984236783E-9 
+PS=839.999984236783E-9 M=1 
M83 2 NCK 4 0  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M84 4 CKDIV 0 0  TSMC25DN  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M85 3 IN 5 0  TSMC25DN  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M86 5 2 0 0  TSMC25DN  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M87 CKDIV 3 0 0  TSMC25DN  L=239.99999143598E-9 W=1.4400000054593E-6 
+AD=864.000006522286E-15 AS=864.000006522286E-15 PD=2.64000004790432E-6 
+PS=2.64000004790432E-6 M=1    
   
.ends   
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dN" NMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc25dP" PMOS 
   
* INCLUDE FILES
   
   
   
   
.END
