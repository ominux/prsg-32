blah

vCLK CLK 0 pulse(0 2.5V 0.5ns 150ps 150ps 0.350ns 1ns )
vVDD VDD! 0 DC 2.5V
vGND GND! 0 DC 0
vRSTIN RSTIN 0 pulse(2.5 0 3.5ns 100ps 100ps 4ns 80ns )
.OPTION list post=2   
.tran 0.01p 80n
.measure tran avgpwr AVG power from=0ns to 80ns
 
.lib 'models25.txt' TT	
   
C85 0 56  26.5392E-18 M=1.0 
C86 0 55  26.5391999999999E-18 M=1.0 
C87 0 23  40.5072000000001E-18 M=1.0 
C88 0 20  46.0943999999999E-18 M=1.0 
C89 0 17  111.744E-18 M=1.0 
C90 0 15  30.3804E-18 M=1.0 
C91 0 12  34.9200000000001E-18 M=1.0 
C92 0 11  36.3168000000002E-18 M=1.0 
C93 0 10  114.5376E-18 M=1.0 
C94 0 9  78.2208E-18 M=1.0 
C95 0 7  114.5376E-18 M=1.0 
C96 0 6  36.3168E-18 M=1.0 
C97 0 5  78.2208E-18 M=1.0 
C98 0 4  34.9200000000001E-18 M=1.0 
C99 0 RST  157.8384E-18 M=1.0 
C100 VDD! 56  47.4912000000001E-18 M=1.0 
C101 VDD! 55  47.4911999999999E-18 M=1.0 
C102 VDD! 26  25.1424E-18 M=1.0 
C103 VDD! 20  23.7455999999999E-18 M=1.0 
C104 VDD! 17  90.792E-18 M=1.0 
C105 VDD! 14  50.2848E-18 M=1.0 
C106 VDD! 13  34.92E-18 M=1.0 
C107 VDD! 12  33.5232E-18 M=1.0 
C108 VDD! 11  34.9199999999999E-18 M=1.0 
C109 VDD! 10  50.2848E-18 M=1.0 
C110 VDD! 9  34.92E-18 M=1.0 
C111 VDD! 8  34.92E-18 M=1.0 
C112 VDD! 7  50.2848E-18 M=1.0 
C113 VDD! 6  34.92E-18 M=1.0 
C114 VDD! 5  34.9199999999999E-18 M=1.0 
C115 VDD! 4  33.5231999999999E-18 M=1.0 
C116 VDD! Q3N  72.6336000000001E-18 M=1.0 
C117 Q6 0  32.1264E-18 M=1.0 
C118 Q6 VDD!  29.3328E-18 M=1.0 
C119 Q5 0  32.1264E-18 M=1.0 
C120 Q5 VDD!  29.3328E-18 M=1.0 
C121 Q2 0  27.936E-18 M=1.0 
C122 Q2 VDD!  43.3007999999999E-18 M=1.0 
C123 CLK 0  194.1552E-18 M=1.0 
C124 NRST 0  76.4747999999999E-18 M=1.0 
C125 NRST VDD!  198.6948E-18 M=1.0 
C126 P4P 0  67.0464E-18 M=1.0 
C127 P4N VDD!  36.3168E-18 M=1.0 
C128 Q7N 0  76.824E-18 M=1.0 
C129 Q7N VDD!  100.5696E-18 M=1.0 
C130 PHN 0  42.6023999999998E-18 M=1.0 
C131 PHI 0  44.6976000000001E-18 M=1.0 
C132 PHI VDD!  33.5232E-18 M=1.0 
C133 P3P 0  148.0608E-18 M=1.0 
C134 P3P VDD!  32.1264E-18 M=1.0 
C135 P3N VDD!  108.9504E-18 M=1.0 
C136 P2P 0  67.0464E-18 M=1.0 
C137 P2P VDD!  32.1264E-18 M=1.0 
C138 P2N VDD!  36.3168E-18 M=1.0 
C139 P1P 0  148.0608E-18 M=1.0 
C140 P1P VDD!  32.1264E-18 M=1.0 
C141 P1N VDD!  108.9504E-18 M=1.0 
C142 Q4N 0  57.2688000000001E-18 M=1.0 
C143 Q4N VDD!  75.4271999999999E-18 M=1.0 
C144 20 21  89.4432E-18 M=1.0 
C145 0 56  51.2496E-18 M=1.0 
C146 0 55  51.2496E-18 M=1.0 
C147 0 21  129.7416E-18 M=1.0 
C148 0 20  125.328E-18 M=1.0 
C149 0 17  233.6568E-18 M=1.0 
C150 0 14  181.3008E-18 M=1.0 
C151 0 13  51.2496E-18 M=1.0 
C152 0 12  157.068E-18 M=1.0 
C153 0 11  133.3584E-18 M=1.0 
C154 0 9  407.9616E-18 M=1.0 
C155 0 8  51.2496E-18 M=1.0 
C156 0 7  135.5952E-18 M=1.0 
C157 0 6  133.3584E-18 M=1.0 
C158 0 5  407.9616E-18 M=1.0 
C159 0 4  157.068E-18 M=1.0 
C160 0 3  149.9424E-18 M=1.0 
C161 0 Q3N  162.624E-18 M=1.0 
C162 0 RST  557.4696E-18 M=1.0 
C163 VDD! 56  144.3504E-18 M=1.0 
C164 VDD! 55  105.3072E-18 M=1.0 
C165 VDD! 23  119.3328E-18 M=1.0 
C166 VDD! 21  137.4624E-18 M=1.0 
C167 VDD! 20  51.2496E-18 M=1.0 
C168 VDD! 17  86.5584E-18 M=1.0 
C169 VDD! 14  126.4464E-18 M=1.0 
C170 VDD! 13  244.6128E-18 M=1.0 
C171 VDD! 12  142.1856E-18 M=1.0 
C172 VDD! 11  151.0368E-18 M=1.0 
C173 VDD! 10  144.0528E-18 M=1.0 
C174 VDD! 9  81.8592E-18 M=1.0 
C175 VDD! 8  244.6128E-18 M=1.0 
C176 VDD! 7  126.4464E-18 M=1.0 
C177 VDD! 6  151.0368E-18 M=1.0 
C178 VDD! 5  81.8592000000001E-18 M=1.0 
C179 VDD! Q3N  123.7344E-18 M=1.0 
C180 Q6 0  101.1552E-18 M=1.0 
C181 Q6 VDD!  141.0912E-18 M=1.0 
C182 Q5 VDD!  141.0912E-18 M=1.0 
C183 Q2 0  99.204E-18 M=1.0 
C184 Q2 VDD!  108.852E-18 M=1.0 
C185 OUT13 0  51.2496E-18 M=1.0 
C186 OUT13 VDD!  51.2496E-18 M=1.0 
C187 CLK 21  126.672E-18 M=1.0 
C188 P4N VDD!  104.1768E-18 M=1.0 
C189 PHN 0  125.1144E-18 M=1.0 
C190 PHI 0  130.6344E-18 M=1.0 
C191 PHI VDD!  81.0264E-18 M=1.0 
C192 P3P 7  89.4432E-18 M=1.0 
C193 P3P VDD!  85.6776E-18 M=1.0 
C194 P3N VDD!  230.9208E-18 M=1.0 
C195 P3N Q7N  232.9152E-18 M=1.0 
C196 P2P 10  89.4432E-18 M=1.0 
C197 P2P 0  126.6672E-18 M=1.0 
C198 P2P VDD!  90.216E-18 M=1.0 
C199 P2N 0  91.7568E-18 M=1.0 
C200 P2N VDD!  104.1768E-18 M=1.0 
C201 P1P 14  89.4432E-18 M=1.0 
C202 P1P 0  330.696E-18 M=1.0 
C203 P1P VDD!  102.9216E-18 M=1.0 
C204 P1N 0  66.132E-18 M=1.0 
C205 P1N VDD!  244.1496E-18 M=1.0 
C206 Q4N 0  146.3496E-18 M=1.0 
C207 Q4N VDD!  148.2408E-18 M=1.0 
C208 OUTGATE 0  147.1584E-18 M=1.0 
C209 OUTGATE VDD!  166.9776E-18 M=1.0 
C210 55 56  135.9888E-18 M=1.0 
C211 12 13  79.6752E-18 M=1.0 
C212 10 16  51.8688E-18 M=1.0 
C213 9 12  254.9436E-18 M=1.0 
C214 8 11  81.1584E-18 M=1.0 
C215 7 10  51.8688E-18 M=1.0 
C216 6 13  81.1584E-18 M=1.0 
C217 6 12  131.544E-18 M=1.0 
C218 4 11  131.544E-18 M=1.0 
C219 4 8  79.6752E-18 M=1.0 
C220 4 5  254.9436E-18 M=1.0 
C221 3 10  103.7376E-18 M=1.0 
C222 0 56  146.1984E-18 M=1.0 
C223 0 55  146.1984E-18 M=1.0 
C224 0 23  51.8688E-18 M=1.0 
C225 0 20  146.1984E-18 M=1.0 
C226 0 13  94.3296E-18 M=1.0 
C227 0 12  566.3568E-18 M=1.0 
C228 0 11  240.528E-18 M=1.0 
C229 0 10  211.0344E-18 M=1.0 
C230 0 9  292.3968E-18 M=1.0 
C231 0 8  94.3296E-18 M=1.0 
C232 0 6  188.6592E-18 M=1.0 
C233 0 5  292.3968E-18 M=1.0 
C234 0 4  472.0272E-18 M=1.0 
C235 0 Q3N  146.4864E-18 M=1.0 
C236 VDD! 56  173.7792E-18 M=1.0 
C237 VDD! 55  194.2416E-18 M=1.0 
C238 VDD! 20  133.0272E-18 M=1.0 
C239 VDD! 12  366.1812E-18 M=1.0 
C240 VDD! 11  53.2728E-18 M=1.0 
C241 VDD! 9  94.6176E-18 M=1.0 
C242 VDD! 6  53.2728E-18 M=1.0 
C243 VDD! 5  94.6176E-18 M=1.0 
C244 VDD! Q3N  198.3552E-18 M=1.0 
C245 VDD! 0  321.228E-18 M=1.0 
C246 Q6 0  146.1984E-18 M=1.0 
C247 Q6 VDD!  146.4864E-18 M=1.0 
C248 Q5 VDD!  146.4864E-18 M=1.0 
C249 Q2 12  51.8688E-18 M=1.0 
C250 Q2 0  146.4864E-18 M=1.0 
C251 Q2 VDD!  51.8688E-18 M=1.0 
C252 Q1 VDD!  94.6176E-18 M=1.0 
C253 OUT13 0  94.9056E-18 M=1.0 
C254 CLK 0  51.8688E-18 M=1.0 
C255 CLK VDD!  103.7376E-18 M=1.0 
C256 NRST 58  93.7536E-18 M=1.0 
C257 NRST RST  105.168E-18 M=1.0 
C258 NRST 0  421.38E-18 M=1.0 
C259 NRST VDD!  281.7048E-18 M=1.0 
C260 P4N VDD!  732.1536E-18 M=1.0 
C261 Q7N P4N  51.8688E-18 M=1.0 
C262 P3P 0  51.8688E-18 M=1.0 
C263 P3N VDD!  103.7376E-18 M=1.0 
C264 P2P 0  863.7624E-18 M=1.0 
C265 P2P VDD!  44.2944E-18 M=1.0 
C266 P2P P3P  421.7784E-18 M=1.0 
C267 P2N 0  372.7224E-18 M=1.0 
C268 P2N VDD!  708.912E-18 M=1.0 
C269 P2N Q7N  36.2592E-18 M=1.0 
C270 P2N P3P  79.6752E-18 M=1.0 
C271 P2N P3N  161.4816E-18 M=1.0 
C272 P1P 0  103.7376E-18 M=1.0 
C273 P1N VDD!  103.7376E-18 M=1.0 
C274 P1N P4N  107.2992E-18 M=1.0 
C275 P1N P2P  228.144E-18 M=1.0 
C276 Q4N 12  51.8688E-18 M=1.0 
C277 Q4N 0  198.3552E-18 M=1.0 
C278 Q4N VDD!  94.6176E-18 M=1.0 
C279 OUTGATE 0  94.3296E-18 M=1.0 
C280 20 22  173.808E-18 M=1.0 
C281 14 17  90.648E-18 M=1.0 
C282 10 14  73.296E-18 M=1.0 
C283 7 14  36.864E-18 M=1.0 
C284 3 10  95.04E-18 M=1.0 
C285 0 17  118.77E-18 M=1.0 
C286 0 14  966.5784E-18 M=1.0 
C287 0 10  77.3832E-18 M=1.0 
C288 0 Q3N  284.5728E-18 M=1.0 
C289 0 RST  515.6664E-18 M=1.0 
C290 VDD! 17  144.066E-18 M=1.0 
C291 VDD! 16  73.728E-18 M=1.0 
C292 VDD! 10  99.3312E-18 M=1.0 
C293 VDD! 7  98.6832E-18 M=1.0 
C294 VDD! RST  480.4752E-18 M=1.0 
C295 Q6 RST  176.112E-18 M=1.0 
C296 Q6 0  199.7208E-18 M=1.0 
C297 Q6 VDD!  90.168E-18 M=1.0 
C298 Q5 RST  176.112E-18 M=1.0 
C299 Q2 0  576.8604E-18 M=1.0 
C300 Q2 VDD!  310.7676E-18 M=1.0 
C301 CLK 22  36.864E-18 M=1.0 
C302 NRST Q3N  222.192E-18 M=1.0 
C303 NRST 0  1.2911712E-15 M=1.0 
C304 NRST VDD!  963.066E-18 M=1.0 
C305 P4P RST  75.4848E-18 M=1.0 
C306 P4N RST  75.4848E-18 M=1.0 
C307 Q7N NRST  102.288E-18 M=1.0 
C308 PHI 9  420.66E-18 M=1.0 
C309 PHI 0  777.0888E-18 M=1.0 
C310 P2P RST  75.4848E-18 M=1.0 
C311 P2P 0  119.238E-18 M=1.0 
C312 P2P VDD!  89.7936E-18 M=1.0 
C313 P2P Q6  75.4848E-18 M=1.0 
C314 P2N RST  75.4848E-18 M=1.0 
C315 P2N P2P  53.784E-18 M=1.0 
C316 P1P 0  1.2988728E-15 M=1.0 
C317 P1P P3P  53.784E-18 M=1.0 
C318 P1P P2P  75.4848E-18 M=1.0 
C319 P1P P2N  75.4848E-18 M=1.0 
C320 Q4N 0  315.1872E-18 M=1.0 
C321 Q4N NRST  222.192E-18 M=1.0 
C322 22 23  79.8048E-18 M=1.0 
C323 20 23  135.5304E-18 M=1.0 
C324 7 14  79.8048E-18 M=1.0 
C325 7 10  291.864E-18 M=1.0 
C326 3 10  217.404E-18 M=1.0 
C327 0 23  106.6032E-18 M=1.0 
C328 0 16  177.3216E-18 M=1.0 
C329 0 10  242.2032E-18 M=1.0 
C330 0 7  179.5488E-18 M=1.0 
C331 VDD! 23  896.6628E-18 M=1.0 
C332 VDD! 16  97.4592E-18 M=1.0 
C333 VDD! 7  29.4048E-18 M=1.0 
C334 VDD! 0  4.40424E-15 M=1.0 
C335 CLK 23  98.5032E-18 M=1.0 
C336 CLK 14  50.2752E-18 M=1.0 
C337 CLK 10  72.1272E-18 M=1.0 
C338 CLK 7  50.2752E-18 M=1.0 
C339 CLK 0  260.424E-18 M=1.0 
C340 PHI VDD!  108.048E-18 M=1.0 
C341 P3P Q3N  79.8048E-18 M=1.0 
C342 P3P RST  79.8048E-18 M=1.0 
C343 P3N RST  79.8048E-18 M=1.0 
C344 P3N VDD!  551.844E-18 M=1.0 
C345 P3N NRST  79.8048E-18 M=1.0 
C346 P3N P4N  637.146E-18 M=1.0 
C347 P3N Q7N  23.8464E-18 M=1.0 
C348 P1P RST  149.8128E-18 M=1.0 
C349 P1P 0  1.432926E-15 M=1.0 
C350 P1P Q6  79.8048E-18 M=1.0 
C351 P1P NRST  252.2712E-18 M=1.0 
C352 P1P Q7N  171.72E-18 M=1.0 
C353 P1P P2P  378.864E-18 M=1.0 
C354 P1N RST  79.8048E-18 M=1.0 
C355 P1N NRST  79.8048E-18 M=1.0 
C356 P1N P2P  79.8048E-18 M=1.0 
C357 P1N P2N  790.7328E-18 M=1.0 
C358 P1N P1P  79.8048E-18 M=1.0 
C359 Q4N P1P  79.8048E-18 M=1.0 
C360 OUTGATE 11  147.6192E-18 M=1.0 
C361 OUTGATE 5  55.0908E-18 M=1.0 
C362 OUTGATE 4  618.4836E-18 M=1.0 
C363 OUTGATE OUT13  42.9264E-18 M=1.0 
C364 16 17  54.0432E-18 M=1.0 
C365 14 17  112.0152E-18 M=1.0 
C366 14 16  76.1328E-18 M=1.0 
C367 10 17  129.8304E-18 M=1.0 
C368 10 16  41.5296E-18 M=1.0 
C369 7 17  541.1136E-18 M=1.0 
C370 7 16  65.4012E-18 M=1.0 
C371 0 17  276.5088E-18 M=1.0 
C372 0 16  1.1500032E-15 M=1.0 
C373 0 15  71.3124E-18 M=1.0 
C374 0 14  46.1808E-18 M=1.0 
C375 0 10  46.1808E-18 M=1.0 
C376 0 7  46.1808E-18 M=1.0 
C377 VDD! 17  141.0048E-18 M=1.0 
C378 VDD! 16  756.0516E-18 M=1.0 
C379 VDD! 14  38.1024E-18 M=1.0 
C380 VDD! 13  103.248E-18 M=1.0 
C381 VDD! 12  63.6768E-18 M=1.0 
C382 VDD! 11  233.5296E-18 M=1.0 
C383 VDD! 10  46.1808E-18 M=1.0 
C384 VDD! 9  46.1808E-18 M=1.0 
C385 VDD! 8  103.248E-18 M=1.0 
C386 VDD! 7  30.5424E-18 M=1.0 
C387 VDD! 6  233.5296E-18 M=1.0 
C388 VDD! 5  46.1808E-18 M=1.0 
C389 VDD! 4  63.6768E-18 M=1.0 
C390 VDD! RST  20.7648E-18 M=1.0 
C391 VDD! 0  1.6477716E-15 M=1.0 
C392 CLK 0  613.8144E-18 M=1.0 
C393 NRST Q3N  66.432E-18 M=1.0 
C394 NRST 0  136.4652E-18 M=1.0 
C395 NRST VDD!  716.0616E-18 M=1.0 
C396 Q7N VDD!  76.488E-18 M=1.0 
C397 P3P 0  245.484E-18 M=1.0 
C398 P3P VDD!  320.694E-18 M=1.0 
C399 P2P 0  282.5544E-18 M=1.0 
C400 P2P VDD!  94.4496E-18 M=1.0 
C401 P2N 0  45.7104E-18 M=1.0 
C402 P2N VDD!  28.4328E-18 M=1.0 
C403 P1P 0  348.264E-18 M=1.0 
C404 P1P VDD!  499.3224E-18 M=1.0 
C405 P1N 0  154.4304E-18 M=1.0 
C406 P1N VDD!  419.3568E-18 M=1.0 
C407 Q4N 0  97.8048E-18 M=1.0 
C408 Q4N VDD!  142.7328E-18 M=1.0 
C409 Q4N Q2  210.528E-18 M=1.0 
C410 Q4N NRST  66.432E-18 M=1.0 
C411 0 14  114.5376E-18 M=1.0 
C412 0 3  114.5376E-18 M=1.0 
C413 0 1  40.5072E-18 M=1.0 
C414 VDD! 3  50.2848E-18 M=1.0 
C415 OUT 0  34.92E-18 M=1.0 
C416 OUT VDD!  26.5392E-18 M=1.0 
C417 P4P VDD!  32.1264E-18 M=1.0 
C418 0 16  145.8384E-18 M=1.0 
C419 0 10  157.6752E-18 M=1.0 
C420 0 2  47.532E-18 M=1.0 
C421 0 1  152.6304E-18 M=1.0 
C422 VDD! 3  152.3088E-18 M=1.0 
C423 VDD! 1  87.6528E-18 M=1.0 
C424 VDD! 0  417.4872E-18 M=1.0 
C425 Q5 0  101.1552E-18 M=1.0 
C426 P4P 3  89.4432E-18 M=1.0 
C427 P4P 0  165.5328E-18 M=1.0 
C428 P4P VDD!  85.6776E-18 M=1.0 
C429 P4N 0  87.6288E-18 M=1.0 
C430 Q7N 0  187.9392E-18 M=1.0 
C431 Q7N VDD!  119.0352E-18 M=1.0 
C432 P3P 0  918.756E-18 M=1.0 
C433 P3N 0  66.132E-18 M=1.0 
C434 3 16  51.8688E-18 M=1.0 
C435 3 14  145.6224E-18 M=1.0 
C436 0 3  410.5608E-18 M=1.0 
C437 Q5 0  146.1984E-18 M=1.0 
C438 P4P 0  812.9088E-18 M=1.0 
C439 P4N 0  449.3736E-18 M=1.0 
C440 Q7N 0  389.214E-18 M=1.0 
C441 Q7N VDD!  325.8168E-18 M=1.0 
C442 Q7N OUT  642.4548E-18 M=1.0 
C443 Q7N CLK  51.8688E-18 M=1.0 
C444 Q7N P4P  93.7536E-18 M=1.0 
C445 P3P P4N  79.6752E-18 M=1.0 
C446 P3N P4N  91.8888E-18 M=1.0 
C447 P1P P4P  93.7536E-18 M=1.0 
C448 VDD! 3  110.1168E-18 M=1.0 
C449 VDD! 0  2.7493956E-15 M=1.0 
C450 Q5 0  347.8608E-18 M=1.0 
C451 Q5 VDD!  90.168E-18 M=1.0 
C452 CLK 1  209.826E-18 M=1.0 
C453 CLK 0  493.1352E-18 M=1.0 
C454 CLK VDD!  145.7532E-18 M=1.0 
C455 P4P Q5  75.4848E-18 M=1.0 
C456 Q7N CLK  75.4848E-18 M=1.0 
C457 P1P VDD!  44.382E-18 M=1.0 
C458 P1P P4P  167.3808E-18 M=1.0 
C459 P1P P4N  134.5608E-18 M=1.0 
C460 P1P Q7N  53.784E-18 M=1.0 
C461 10 14  117.9216E-18 M=1.0 
C462 VDD! 3  29.4048E-18 M=1.0 
C463 VDD! 1  53.9496E-18 M=1.0 
C464 OUT VDD!  105.9348E-18 M=1.0 
C465 CLK 57  50.2752E-18 M=1.0 
C466 CLK 3  72.1272E-18 M=1.0 
C467 CLK 2  132.5052E-18 M=1.0 
C468 P4P VDD!  50.7648E-18 M=1.0 
C469 Q7N VDD!  96.7104E-18 M=1.0 
C470 P3P 0  497.9088E-18 M=1.0 
C471 P3P Q5  79.8048E-18 M=1.0 
C472 P3P P4P  342.684E-18 M=1.0 
C473 P3N 0  188.9712E-18 M=1.0 
C474 P1P VDD!  448.8936E-18 M=1.0 
C475 P1P Q5  79.8048E-18 M=1.0 
C476 P1P P3P  79.8048E-18 M=1.0 
C477 P1P P3N  142.1208E-18 M=1.0 
C478 0 3  46.1808E-18 M=1.0 
C479 0 2  43.2648E-18 M=1.0 
C480 0 1  80.2944E-18 M=1.0 
C481 VDD! 3  22.8528E-18 M=1.0 
C482 Q5 0  56.1888E-18 M=1.0 
C483 P4P 0  136.104E-18 M=1.0 
C484 P4P VDD!  46.1808E-18 M=1.0 
C485 P4N 0  129.276E-18 M=1.0 
C486 P4N VDD!  57.3048E-18 M=1.0 
C487 Q7N 0  206.6544E-18 M=1.0 
C488 P3N 0  142.5828E-18 M=1.0 
C489 P3N VDD!  281.7696E-18 M=1.0 
C490 0 Q3N  60.0624E-18 M=1.0 
C491 Q1 0  27.936E-18 M=1.0 
C492 Q1 VDD!  43.3008E-18 M=1.0 
C493 PHN VDD!  35.6184E-18 M=1.0 
C494 OUTGATE 0  33.5232E-18 M=1.0 
C495 OUTGATE VDD!  32.1263999999999E-18 M=1.0 
C496 VDD! 4  142.1856E-18 M=1.0 
C497 Q1 0  531.3744E-18 M=1.0 
C498 Q1 VDD!  200.2992E-18 M=1.0 
C499 OUT 0  1.3233744E-15 M=1.0 
C500 OUT VDD!  233.8128E-18 M=1.0 
C501 PHN VDD!  97.0152E-18 M=1.0 
C502 OUT24F 0  51.2496E-18 M=1.0 
C503 OUT24F VDD!  51.2496E-18 M=1.0 
C504 Q3N 4  51.8688E-18 M=1.0 
C505 VDD! 4  366.1812E-18 M=1.0 
C506 Q1 4  51.8688E-18 M=1.0 
C507 OUT 0  478.6968E-18 M=1.0 
C508 PHN 0  3.2199696E-15 M=1.0 
C509 PHN VDD!  625.0632E-18 M=1.0 
C510 PHN Q1  637.4016E-18 M=1.0 
C511 PHN OUT  57.3696E-18 M=1.0 
C512 OUTGATE PHN  51.8688E-18 M=1.0 
C513 VDD! 4  63.6696E-18 M=1.0 
C514 Q1 VDD!  36.864E-18 M=1.0 
C515 OUT 0  163.6188E-18 M=1.0 
C516 OUT VDD!  231.5232E-18 M=1.0 
C517 PHN 0  138.3264E-18 M=1.0 
C518 PHN VDD!  75.4848E-18 M=1.0 
C519 PHI Q1  97.74E-18 M=1.0 
C520 PHI PHN  285.5328E-18 M=1.0 
C521 P3P 0  36.864E-18 M=1.0 
C522 OUTGATE VDD!  36.864E-18 M=1.0 
C523 OUTGATE OUT  36.864E-18 M=1.0 
C524 P3P VDD!  837.9984E-18 M=1.0 
C525 P3P Q1  31.6584E-18 M=1.0 
C526 P3P NRST  420.528E-18 M=1.0 
C527 P3P PHN  155.952E-18 M=1.0 
C528 P3N Q1  183.7008E-18 M=1.0 
C529 P1P OUT  277.9524E-18 M=1.0 
C530 P1P PHN  230.256E-18 M=1.0 
C531 P1N 0  122.9328E-18 M=1.0 
C532 P1N VDD!  973.8576E-18 M=1.0 
C533 P1N Q1  25.1376E-18 M=1.0 
C534 P1N PHN  209.0016E-18 M=1.0 
C535 P1N PHI  50.7504E-18 M=1.0 
C536 P1N P3N  43.584E-18 M=1.0 
C537 OUTGATE 0  523.6416E-18 M=1.0 
C538 OUTGATE VDD!  563.8896E-18 M=1.0 
C539 OUTGATE Q1  115.6776E-18 M=1.0 
C540 OUTGATE OUT  42.9264E-18 M=1.0 
C541 OUTGATE PHN  235.332E-18 M=1.0 
C542 OUTGATE PHI  275.2128E-18 M=1.0 
C543 0 Q3N  276.9696E-18 M=1.0 
C544 VDD! Q3N  234.0288E-18 M=1.0 
C545 Q1 Q3N  50.22E-18 M=1.0 
C546 PHN Q3N  98.736E-18 M=1.0 
C547 PHI Q3N  143.136E-18 M=1.0 
C548 P3N Q3N  115.5936E-18 M=1.0 
C549 P1N Q3N  115.5936E-18 M=1.0 
C550 0 21  55.8720000000001E-18 M=1.0 
C551 0 16  92.1888000000001E-18 M=1.0 
C552 VDD! 21  23.7456000000001E-18 M=1.0 
C553 VDD! 16  110.3472E-18 M=1.0 
C554 VDD! 15  40.8564E-18 M=1.0 
C555 VDD! RST  34.92E-18 M=1.0 
C556 CLK VDD!  257.0112E-18 M=1.0 
C557 RSTIN VDD!  148.0608E-18 M=1.0 
C558 RST 21  89.4432E-18 M=1.0 
C559 0 26  483.9912E-18 M=1.0 
C560 0 23  92.8752E-18 M=1.0 
C561 0 15  83.9232E-18 M=1.0 
C562 VDD! 26  51.2496E-18 M=1.0 
C563 VDD! 22  51.2496E-18 M=1.0 
C564 VDD! 16  203.0832E-18 M=1.0 
C565 VDD! 15  94.9392E-18 M=1.0 
C566 VDD! RST  195.1128E-18 M=1.0 
C567 CLK 0  253.62E-18 M=1.0 
C568 CLK VDD!  793.9392E-18 M=1.0 
C569 NRST 0  395.5488E-18 M=1.0 
C570 NRST VDD!  174.1872E-18 M=1.0 
C571 RST 21  79.6752E-18 M=1.0 
C572 0 21  237.8112E-18 M=1.0 
C573 0 RST  160.2768E-18 M=1.0 
C574 VDD! 26  146.4864E-18 M=1.0 
C575 VDD! 21  214.1856E-18 M=1.0 
C576 VDD! RST  159.7656E-18 M=1.0 
C577 RSTIN 0  51.8688E-18 M=1.0 
C578 RSTIN VDD!  937.2612E-18 M=1.0 
C579 21 22  321.0504E-18 M=1.0 
C580 15 17  90.648E-18 M=1.0 
C581 15 16  90.648E-18 M=1.0 
C582 RST 22  73.044E-18 M=1.0 
C583 0 22  870.4296E-18 M=1.0 
C584 0 15  265.7304E-18 M=1.0 
C585 VDD! 15  269.3808E-18 M=1.0 
C586 CLK 15  73.728E-18 M=1.0 
C587 NRST 22  90.648E-18 M=1.0 
C588 15 16  79.8048E-18 M=1.0 
C589 CLK 15  243.1368E-18 M=1.0 
C590 CLK VDD!  1.1983104E-15 M=1.0 
C591 0 23  115.5936E-18 M=1.0 
C592 0 22  66.432E-18 M=1.0 
C593 0 21  45.9588E-18 M=1.0 
C594 0 RST  129.8088E-18 M=1.0 
C595 VDD! 23  50.5728E-18 M=1.0 
C596 VDD! 15  61.4448E-18 M=1.0 
C597 CLK VDD!  207.9552E-18 M=1.0 
C598 0 27  34.9200000000001E-18 M=1.0 
C599 0 26  92.1887999999999E-18 M=1.0 
C600 0 25  34.9200000000001E-18 M=1.0 
C601 0 22  54.4751999999999E-18 M=1.0 
C602 0 19  122.22E-18 M=1.0 
C603 0 18  37.7136E-18 M=1.0 
C604 VDD! 27  33.5232E-18 M=1.0 
C605 VDD! 25  26.5392E-18 M=1.0 
C606 VDD! 24  34.92E-18 M=1.0 
C607 VDD! 19  67.0463999999999E-18 M=1.0 
C608 VDD! 18  34.9200000000001E-18 M=1.0 
C609 RSTIN 0  54.4752E-18 M=1.0 
C610 18 19  89.4432E-18 M=1.0 
C611 0 27  92.5896E-18 M=1.0 
C612 0 25  161.0352E-18 M=1.0 
C613 0 24  51.2496E-18 M=1.0 
C614 0 22  139.9848E-18 M=1.0 
C615 0 19  146.1528E-18 M=1.0 
C616 0 18  183.0792E-18 M=1.0 
C617 VDD! 27  76.6128E-18 M=1.0 
C618 VDD! 25  174.0864E-18 M=1.0 
C619 VDD! 24  193.6608E-18 M=1.0 
C620 VDD! 19  103.5816E-18 M=1.0 
C621 VDD! 18  224.472E-18 M=1.0 
C622 RSTIN VDD!  731.4408E-18 M=1.0 
C623 25 27  131.544E-18 M=1.0 
C624 24 25  51.8688E-18 M=1.0 
C625 18 19  131.544E-18 M=1.0 
C626 0 27  250.0704E-18 M=1.0 
C627 0 26  291.0432E-18 M=1.0 
C628 0 25  158.8608E-18 M=1.0 
C629 0 22  51.8688E-18 M=1.0 
C630 0 19  418.8288E-18 M=1.0 
C631 0 18  247.1676E-18 M=1.0 
C632 VDD! 27  118.4832E-18 M=1.0 
C633 VDD! 25  53.2728E-18 M=1.0 
C634 VDD! 24  147.3504E-18 M=1.0 
C635 VDD! 19  211.6344E-18 M=1.0 
C636 VDD! 18  241.536E-18 M=1.0 
C637 RSTIN 25  81.1584E-18 M=1.0 
C638 RSTIN 24  51.8688E-18 M=1.0 
C639 19 22  484.9644E-18 M=1.0 
C640 18 22  116.82E-18 M=1.0 
C641 VDD! 22  66.432E-18 M=1.0 
C642 VDD! 19  25.1376E-18 M=1.0 
C643 VDD! 18  131.3928E-18 M=1.0 
M644 OUT OUTGATE VDD! VDD!  pmos  L=239.99999143598E-9 
+W=2.15999989450211E-6 AD=1.29599998267838E-12 AS=1.29599998267838E-12 
+PD=3.35999993694713E-6 PS=3.35999993694713E-6 M=1 
M645 P1P 14 VDD! VDD!  pmos  L=239.99999143598E-9 W=600.000021222513E-9 
+AD=417.600009476951E-15 AS=251.999999643579E-15 PD=2.04000002668181E-6 
+PS=779.999993483216E-9 M=1 
M646 VDD! 10 P2P VDD!  pmos  L=239.99999143598E-9 W=600.000021222513E-9 
+AD=251.999999643579E-15 AS=417.600009476951E-15 PD=779.999993483216E-9 
+PS=2.04000002668181E-6 M=1 
M647 P3P 7 VDD! VDD!  pmos  L=239.99999143598E-9 W=600.000021222513E-9 
+AD=417.600009476951E-15 AS=251.999999643579E-15 PD=2.04000002668181E-6 
+PS=779.999993483216E-9 M=1 
M648 VDD! 3 P4P VDD!  pmos  L=239.99999143598E-9 W=600.000021222513E-9 
+AD=251.999999643579E-15 AS=417.600009476951E-15 PD=779.999993483216E-9 
+PS=2.04000002668181E-6 M=1 
M649 12 Q4N VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=259.199996535675E-15 PD=1.91999993148784E-6 
+PS=720.000002729648E-9 M=1 
M650 OUTGATE PHI OUT13 VDD!  pmos  L=239.99999143598E-9 
+W=720.000002729648E-9 AD=432.000003261143E-15 AS=259.199996535675E-15 
+PD=1.91999993148784E-6 PS=720.000002729648E-9 M=1 
M651 VDD! Q2 9 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=432.000003261143E-15 PD=720.000002729648E-9 
+PS=1.91999993148784E-6 M=1 
M652 OUT13 11 VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=432.000003261143E-15 PD=720.000002729648E-9 
+PS=1.91999993148784E-6 M=1 
M653 VDD! P1P P1N VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=251.999999643579E-15 AS=432.000003261143E-15 PD=779.999993483216E-9 
+PS=1.91999993148784E-6 M=1 
M654 VDD! 9 13 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=432.000003261143E-15 PD=1.91999993148784E-6 
+PS=1.91999993148784E-6 M=1 
M655 11 4 8 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=432.000003261143E-15 PD=1.91999993148784E-6 
+PS=1.91999993148784E-6 M=1 
M656 P2N P2P VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=251.999999643579E-15 PD=1.91999993148784E-6 
+PS=779.999993483216E-9 M=1 
M657 12 13 6 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=432.000003261143E-15 PD=1.91999993148784E-6 
+PS=1.91999993148784E-6 M=1 
M658 11 8 4 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=432.000003261143E-15 PD=1.91999993148784E-6 
+PS=1.91999993148784E-6 M=1 
M659 13 12 6 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=432.000003261143E-15 PD=1.91999993148784E-6 
+PS=1.91999993148784E-6 M=1 
M660 8 5 VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=432.000003261143E-15 PD=1.91999993148784E-6 
+PS=1.91999993148784E-6 M=1 
M661 VDD! 6 OUT24F VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=259.199996535675E-15 PD=1.91999993148784E-6 
+PS=720.000002729648E-9 M=1 
M662 VDD! P3P P3N VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=251.999999643579E-15 AS=432.000003261143E-15 PD=779.999993483216E-9 
+PS=1.91999993148784E-6 M=1 
M663 5 Q3N VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=259.199996535675E-15 PD=1.91999993148784E-6 
+PS=720.000002729648E-9 M=1 
M664 OUT24F PHN OUTGATE VDD!  pmos  L=239.99999143598E-9 
+W=720.000002729648E-9 AD=259.199996535675E-15 AS=432.000003261143E-15 
+PD=720.000002729648E-9 PS=1.91999993148784E-6 M=1 
M665 VDD! Q1 4 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=432.000003261143E-15 PD=720.000002729648E-9 
+PS=1.91999993148784E-6 M=1 
M666 P4N P4P VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=251.999999643579E-15 PD=1.91999993148784E-6 
+PS=779.999993483216E-9 M=1 
M667 PHI P3N VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=259.199996535675E-15 PD=1.91999993148784E-6 
+PS=720.000002729648E-9 M=1 
M668 VDD! P1N PHN VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=432.000003261143E-15 PD=720.000002729648E-9 
+PS=1.91999993148784E-6 M=1 
M669 Q7N CLK 77 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M670 77 OUT VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M671 18 24 VDD! VDD!  pmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=712.799990473106E-15 AS=647.999991339188E-15 PD=2.40000008489005E-6 
+PS=2.27999998969608E-6 M=1 
M672 18 19 VDD! VDD!  pmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M673 57 CLK 1 VDD!  pmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M674 VDD! CLK 23 VDD!  pmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M675 58 NRST Q6 VDD!  pmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M676 VDD! NRST Q2 VDD!  pmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M677 14 17 VDD! VDD!  pmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M678 VDD! 16 10 VDD!  pmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M679 7 17 VDD! VDD!  pmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M680 VDD! 16 3 VDD!  pmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M681 Q1 NRST VDD! VDD!  pmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M682 Q5 NRST VDD! VDD!  pmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M683 VDD! RSTIN 24 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=432.000003261143E-15 PD=720.000002729648E-9 
+PS=1.91999993148784E-6 M=1 
M684 26 RSTIN VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=259.199996535675E-15 PD=1.91999993148784E-6 
+PS=720.000002729648E-9 M=1 
M685 VDD! 26 56 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=432.000003261143E-15 PD=720.000002729648E-9 
+PS=1.91999993148784E-6 M=1 
M686 55 56 VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=259.199996535675E-15 PD=1.91999993148784E-6 
+PS=720.000002729648E-9 M=1 
M687 VDD! 55 27 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=259.199996535675E-15 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M688 27 RSTIN 25 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=432.000003261143E-15 PD=720.000002729648E-9 
+PS=1.91999993148784E-6 M=1 
M689 RSTIN 27 25 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=432.000003261143E-15 PD=1.91999993148784E-6 
+PS=1.91999993148784E-6 M=1 
M690 24 25 VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=259.199996535675E-15 PD=1.91999993148784E-6 
+PS=720.000002729648E-9 M=1 
M691 22 NRST VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=432.000003261143E-15 PD=1.91999993148784E-6 
+PS=1.91999993148784E-6 M=1 
M692 NRST RST VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=259.199996535675E-15 PD=1.91999993148784E-6 
+PS=720.000002729648E-9 M=1 
M693 VDD! 21 RST VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=432.000003261143E-15 PD=720.000002729648E-9 
+PS=1.91999993148784E-6 M=1 
M694 21 CLK VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=259.199996535675E-15 PD=1.91999993148784E-6 
+PS=720.000002729648E-9 M=1 
M695 VDD! 20 21 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=432.000003261143E-15 PD=720.000002729648E-9 
+PS=1.91999993148784E-6 M=1 
M696 20 CLK 84 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M697 84 19 VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M698 19 18 VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=432.000003261143E-15 PD=1.91999993148784E-6 
+PS=1.91999993148784E-6 M=1 
M699 VDD! 15 17 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=259.199996535675E-15 PD=1.91999993148784E-6 
+PS=720.000002729648E-9 M=1 
M700 17 16 VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=259.199996535675E-15 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M701 VDD! 17 16 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=259.199996535675E-15 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M702 16 CLK VDD! VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=259.199996535675E-15 PD=720.000002729648E-9 
+PS=720.000002729648E-9 M=1 
M703 VDD! CLK 15 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=259.199996535675E-15 AS=432.000003261143E-15 PD=720.000002729648E-9 
+PS=1.91999993148784E-6 M=1 
M704 83 P3N Q6 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M705 VDD! Q6 82 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M706 82 P2N Q4N VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M707 VDD! Q4N 81 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M708 81 P1N Q2 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M709 VDD! Q7N 83 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M710 VDD! Q7N 80 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M711 80 P1N Q5 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M712 VDD! Q5 79 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M713 79 P4N Q3N VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M714 VDD! Q3N 78 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M715 78 P3N Q1 VDD!  pmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M716 OUT OUTGATE 0 0  nmos  L=239.99999143598E-9 W=1.07999994725105E-6 
+AD=647.999991339188E-15 AS=647.999991339188E-15 PD=2.27999998969608E-6 
+PS=2.27999998969608E-6 M=1 
M717 P1P 14 0 0  nmos  L=239.99999143598E-9 W=600.000021222513E-9 
+AD=360.000007235128E-15 AS=201.599994293852E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M718 0 10 P2P 0  nmos  L=239.99999143598E-9 W=600.000021222513E-9 
+AD=201.599994293852E-15 AS=360.000007235128E-15 PD=839.999984236783E-9 
+PS=1.7999999499807E-6 M=1 
M719 P3P 7 0 0  nmos  L=239.99999143598E-9 W=600.000021222513E-9 
+AD=360.000007235128E-15 AS=201.599994293852E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M720 0 3 P4P 0  nmos  L=239.99999143598E-9 W=600.000021222513E-9 
+AD=201.599994293852E-15 AS=360.000007235128E-15 PD=839.999984236783E-9 
+PS=1.7999999499807E-6 M=1 
M721 21 CLK 74 0  nmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=432.000003261143E-15 AS=172.800006725468E-15 PD=1.91999993148784E-6 
+PS=479.999982871959E-9 M=1 
M722 74 20 0 0  nmos  L=239.99999143598E-9 W=720.000002729648E-9 
+AD=172.800006725468E-15 AS=432.000003261143E-15 PD=479.999982871959E-9 
+PS=1.91999993148784E-6 M=1 
M723 18 19 0 0  nmos  L=600.000021222513E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M724 0 CLK 23 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M725 12 Q4N 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=158.399999388749E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M726 0 RST Q4N 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M727 OUTGATE PHN OUT13 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=158.399999388749E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M728 0 Q2 9 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=273.599990319867E-15 PD=839.999984236783E-9 
+PS=1.7999999499807E-6 M=1 
M729 OUT13 11 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=273.599990319867E-15 PD=839.999984236783E-9 
+PS=1.7999999499807E-6 M=1 
M730 14 7 73 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M731 73 17 72 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=86.4000033627341E-15 PD=479.999982871959E-9 
+PS=479.999982871959E-9 M=1 
M732 0 P1P P1N 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=201.599994293852E-15 AS=273.599990319867E-15 PD=839.999984236783E-9 
+PS=1.7999999499807E-6 M=1 
M733 0 9 13 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M734 72 10 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=158.399999388749E-15 PD=479.999982871959E-9 
+PS=839.999984236783E-9 M=1 
M735 11 4 5 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M736 0 7 68 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=86.4000033627341E-15 PD=839.999984236783E-9 
+PS=479.999982871959E-9 M=1 
M737 68 16 67 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=86.4000033627341E-15 PD=479.999982871959E-9 
+PS=479.999982871959E-9 M=1 
M738 12 9 6 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M739 P2N P2P 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=201.599994293852E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M740 11 5 4 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M741 67 3 10 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M742 9 12 6 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M743 8 5 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M744 7 14 66 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M745 66 17 65 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=86.4000033627341E-15 PD=479.999982871959E-9 
+PS=479.999982871959E-9 M=1 
M746 0 6 OUT24F 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=158.399999388749E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M747 65 3 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=158.399999388749E-15 PD=479.999982871959E-9 
+PS=839.999984236783E-9 M=1 
M748 0 P3P P3N 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=201.599994293852E-15 AS=273.599990319867E-15 PD=839.999984236783E-9 
+PS=1.7999999499807E-6 M=1 
M749 5 Q3N 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=158.399999388749E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M750 0 14 64 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=86.4000033627341E-15 PD=839.999984236783E-9 
+PS=479.999982871959E-9 M=1 
M751 OUT24F PHI OUTGATE 0  nmos  L=239.99999143598E-9 
+W=360.000001364824E-9 AD=158.399999388749E-15 AS=273.599990319867E-15 
+PD=839.999984236783E-9 PS=1.7999999499807E-6 M=1 
M752 0 Q1 4 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=273.599990319867E-15 PD=839.999984236783E-9 
+PS=1.7999999499807E-6 M=1 
M753 64 16 60 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=86.4000033627341E-15 PD=479.999982871959E-9 
+PS=479.999982871959E-9 M=1 
M754 P4N P4P 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=201.599994293852E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M755 60 10 3 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M756 Q3N RST 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M757 PHI P1P 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=158.399999388749E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M758 0 P3P PHN 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=273.599990319867E-15 PD=839.999984236783E-9 
+PS=1.7999999499807E-6 M=1 
M759 Q7N 1 59 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M760 0 RST Q7N 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M761 59 OUT 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M762 76 RSTIN 24 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M763 0 25 76 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M764 26 RSTIN 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=158.399999388749E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M765 0 26 56 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=273.599990319867E-15 PD=839.999984236783E-9 
+PS=1.7999999499807E-6 M=1 
M766 55 56 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=158.399999388749E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M767 0 55 27 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=158.399999388749E-15 PD=839.999984236783E-9 
+PS=839.999984236783E-9 M=1 
M768 27 26 25 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=273.599990319867E-15 PD=839.999984236783E-9 
+PS=1.7999999499807E-6 M=1 
M769 26 27 25 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M770 20 23 75 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M771 75 19 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M772 19 18 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M773 18 22 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M774 22 NRST 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
M775 NRST RST 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=158.399999388749E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M776 0 21 RST 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=273.599990319867E-15 PD=839.999984236783E-9 
+PS=1.7999999499807E-6 M=1 
M777 0 CLK 15 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=273.599990319867E-15 PD=839.999984236783E-9 
+PS=1.7999999499807E-6 M=1 
M778 0 15 17 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=158.399999388749E-15 PD=1.7999999499807E-6 
+PS=839.999984236783E-9 M=1 
M779 17 16 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=158.399999388749E-15 PD=839.999984236783E-9 
+PS=839.999984236783E-9 M=1 
M780 0 17 16 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=158.399999388749E-15 PD=839.999984236783E-9 
+PS=839.999984236783E-9 M=1 
M781 16 CLK 0 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=158.399999388749E-15 AS=158.399999388749E-15 PD=839.999984236783E-9 
+PS=839.999984236783E-9 M=1 
M782 0 Q7N 71 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M783 71 P3P Q6 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M784 0 Q6 70 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M785 70 P2P Q4N 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M786 0 Q4N 69 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M787 69 P1P Q2 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M788 61 P3P Q1 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M789 0 Q7N 63 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M790 63 P1P Q5 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M791 0 Q5 62 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M792 62 P4P Q3N 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=86.4000033627341E-15 AS=273.599990319867E-15 PD=479.999982871959E-9 
+PS=1.7999999499807E-6 M=1 
M793 0 Q3N 61 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=86.4000033627341E-15 PD=1.7999999499807E-6 
+PS=479.999982871959E-9 M=1 
M794 2 CLK 1 0  nmos  L=239.99999143598E-9 W=360.000001364824E-9 
+AD=273.599990319867E-15 AS=273.599990319867E-15 PD=1.7999999499807E-6 
+PS=1.7999999499807E-6 M=1 
   
   
   
   

.END
